/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408c80; // 00400014: SLL, REG[17]<=REG[0]<<18;
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdff48; // 00400020: ADDIU, REG[29]<=REG[29]+65352(=0x0000ff48);
      10'h009: data = 32'hafbf00b4; // 00400024: SW, RAM[REG[29]+180]<=REG[31];
      10'h00a: data = 32'hafbe00b0; // 00400028: SW, RAM[REG[29]+176]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h3c020001; // 00400030: LUI
      10'h00d: data = 32'h344286a0; // 00400034: ORI, REG[2]<=REG[2]|0x000086a0;
      10'h00e: data = 32'hafc20010; // 00400038: SW, RAM[REG[30]+16]<=REG[2];
      10'h00f: data = 32'h8fc20010; // 0040003c: LW, REG[2]<=RAM[REG[30]+16];
      10'h010: data = 32'h00000000; // 00400040: SLL, REG[0]<=REG[0]<<0;
      10'h011: data = 32'h00021080; // 00400044: SLL, REG[2]<=REG[2]<<2;
      10'h012: data = 32'h24420007; // 00400048: ADDIU, REG[2]<=REG[2]+7(=0x00000007);
      10'h013: data = 32'h24420007; // 0040004c: ADDIU, REG[2]<=REG[2]+7(=0x00000007);
      10'h014: data = 32'h000210c2; // 00400050: SRL, REG[2]<=REG[2]>>3;
      10'h015: data = 32'h000210c0; // 00400054: SLL, REG[2]<=REG[2]<<3;
      10'h016: data = 32'h03a2e823; // 00400058: SUBU, REG[29]<=REG[29]-REG[2];
      10'h017: data = 32'h27a20010; // 0040005c: ADDIU, REG[2]<=REG[29]+16(=0x00000010);
      10'h018: data = 32'hafc200a8; // 00400060: SW, RAM[REG[30]+168]<=REG[2];
      10'h019: data = 32'h8fc300a8; // 00400064: LW, REG[3]<=RAM[REG[30]+168];
      10'h01a: data = 32'h00000000; // 00400068: SLL, REG[0]<=REG[0]<<0;
      10'h01b: data = 32'h24620007; // 0040006c: ADDIU, REG[2]<=REG[3]+7(=0x00000007);
      10'h01c: data = 32'h000210c2; // 00400070: SRL, REG[2]<=REG[2]>>3;
      10'h01d: data = 32'h000210c0; // 00400074: SLL, REG[2]<=REG[2]<<3;
      10'h01e: data = 32'hafc200a8; // 00400078: SW, RAM[REG[30]+168]<=REG[2];
      10'h01f: data = 32'h8fc200a8; // 0040007c: LW, REG[2]<=RAM[REG[30]+168];
      10'h020: data = 32'h00000000; // 00400080: SLL, REG[0]<=REG[0]<<0;
      10'h021: data = 32'hafc20020; // 00400084: SW, RAM[REG[30]+32]<=REG[2];
      10'h022: data = 32'hafc0001c; // 00400088: SW, RAM[REG[30]+28]<=REG[0];
      10'h023: data = 32'h0810002f; // 0040008c: J, PC<=0x0010002f*4(=0x004000bc);
      10'h024: data = 32'h00000000; // 00400090: SLL, REG[0]<=REG[0]<<0;
      10'h025: data = 32'h8fc2001c; // 00400094: LW, REG[2]<=RAM[REG[30]+28];
      10'h026: data = 32'h8fc30020; // 00400098: LW, REG[3]<=RAM[REG[30]+32];
      10'h027: data = 32'h00021080; // 0040009c: SLL, REG[2]<=REG[2]<<2;
      10'h028: data = 32'h00431821; // 004000a0: ADDU, REG[3]<=REG[2]+REG[3];
      10'h029: data = 32'h24020001; // 004000a4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h02a: data = 32'hac620000; // 004000a8: SW, RAM[REG[3]+0]<=REG[2];
      10'h02b: data = 32'h8fc2001c; // 004000ac: LW, REG[2]<=RAM[REG[30]+28];
      10'h02c: data = 32'h00000000; // 004000b0: SLL, REG[0]<=REG[0]<<0;
      10'h02d: data = 32'h24420001; // 004000b4: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h02e: data = 32'hafc2001c; // 004000b8: SW, RAM[REG[30]+28]<=REG[2];
      10'h02f: data = 32'h8fc2001c; // 004000bc: LW, REG[2]<=RAM[REG[30]+28];
      10'h030: data = 32'h8fc30010; // 004000c0: LW, REG[3]<=RAM[REG[30]+16];
      10'h031: data = 32'h00000000; // 004000c4: SLL, REG[0]<=REG[0]<<0;
      10'h032: data = 32'h0043102b; // 004000c8: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h033: data = 32'h1440fff1; // 004000cc: BNE, PC<=(REG[2] != REG[0])?PC+4+65521*4:PC+4;
      10'h034: data = 32'h00000000; // 004000d0: SLL, REG[0]<=REG[0]<<0;
      10'h035: data = 32'h24020048; // 004000d4: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h036: data = 32'hafc20024; // 004000d8: SW, RAM[REG[30]+36]<=REG[2];
      10'h037: data = 32'h24020045; // 004000dc: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h038: data = 32'hafc20028; // 004000e0: SW, RAM[REG[30]+40]<=REG[2];
      10'h039: data = 32'h2402004c; // 004000e4: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h03a: data = 32'hafc2002c; // 004000e8: SW, RAM[REG[30]+44]<=REG[2];
      10'h03b: data = 32'h2402004c; // 004000ec: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h03c: data = 32'hafc20030; // 004000f0: SW, RAM[REG[30]+48]<=REG[2];
      10'h03d: data = 32'h2402004f; // 004000f4: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h03e: data = 32'hafc20034; // 004000f8: SW, RAM[REG[30]+52]<=REG[2];
      10'h03f: data = 32'h2402000a; // 004000fc: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h040: data = 32'hafc20038; // 00400100: SW, RAM[REG[30]+56]<=REG[2];
      10'h041: data = 32'hafc0003c; // 00400104: SW, RAM[REG[30]+60]<=REG[0];
      10'h042: data = 32'h27c20024; // 00400108: ADDIU, REG[2]<=REG[30]+36(=0x00000024);
      10'h043: data = 32'h00402021; // 0040010c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h044: data = 32'h0c100257; // 00400110: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h045: data = 32'h00000000; // 00400114: SLL, REG[0]<=REG[0]<<0;
      10'h046: data = 32'h2402004e; // 00400118: ADDIU, REG[2]<=REG[0]+78(=0x0000004e);
      10'h047: data = 32'hafc20024; // 0040011c: SW, RAM[REG[30]+36]<=REG[2];
      10'h048: data = 32'h24020055; // 00400120: ADDIU, REG[2]<=REG[0]+85(=0x00000055);
      10'h049: data = 32'hafc20028; // 00400124: SW, RAM[REG[30]+40]<=REG[2];
      10'h04a: data = 32'h2402004d; // 00400128: ADDIU, REG[2]<=REG[0]+77(=0x0000004d);
      10'h04b: data = 32'hafc2002c; // 0040012c: SW, RAM[REG[30]+44]<=REG[2];
      10'h04c: data = 32'h2402003d; // 00400130: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h04d: data = 32'hafc20030; // 00400134: SW, RAM[REG[30]+48]<=REG[2];
      10'h04e: data = 32'hafc00034; // 00400138: SW, RAM[REG[30]+52]<=REG[0];
      10'h04f: data = 32'h27c20024; // 0040013c: ADDIU, REG[2]<=REG[30]+36(=0x00000024);
      10'h050: data = 32'h00402021; // 00400140: ADDU, REG[4]<=REG[2]+REG[0];
      10'h051: data = 32'h0c100257; // 00400144: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h052: data = 32'h00000000; // 00400148: SLL, REG[0]<=REG[0]<<0;
      10'h053: data = 32'h27c20064; // 0040014c: ADDIU, REG[2]<=REG[30]+100(=0x00000064);
      10'h054: data = 32'h00402021; // 00400150: ADDU, REG[4]<=REG[2]+REG[0];
      10'h055: data = 32'h0c100175; // 00400154: JAL, PC<=0x00100175*4(=0x004005d4); REG[31]<=PC+4
      10'h056: data = 32'h00000000; // 00400158: SLL, REG[0]<=REG[0]<<0;
      10'h057: data = 32'h24020045; // 0040015c: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h058: data = 32'hafc20024; // 00400160: SW, RAM[REG[30]+36]<=REG[2];
      10'h059: data = 32'h24020043; // 00400164: ADDIU, REG[2]<=REG[0]+67(=0x00000043);
      10'h05a: data = 32'hafc20028; // 00400168: SW, RAM[REG[30]+40]<=REG[2];
      10'h05b: data = 32'h24020048; // 0040016c: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h05c: data = 32'hafc2002c; // 00400170: SW, RAM[REG[30]+44]<=REG[2];
      10'h05d: data = 32'h2402004f; // 00400174: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h05e: data = 32'hafc20030; // 00400178: SW, RAM[REG[30]+48]<=REG[2];
      10'h05f: data = 32'h24020020; // 0040017c: ADDIU, REG[2]<=REG[0]+32(=0x00000020);
      10'h060: data = 32'hafc20034; // 00400180: SW, RAM[REG[30]+52]<=REG[2];
      10'h061: data = 32'hafc00038; // 00400184: SW, RAM[REG[30]+56]<=REG[0];
      10'h062: data = 32'h27c20024; // 00400188: ADDIU, REG[2]<=REG[30]+36(=0x00000024);
      10'h063: data = 32'h00402021; // 0040018c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h064: data = 32'h0c100257; // 00400190: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h065: data = 32'h00000000; // 00400194: SLL, REG[0]<=REG[0]<<0;
      10'h066: data = 32'h27c20064; // 00400198: ADDIU, REG[2]<=REG[30]+100(=0x00000064);
      10'h067: data = 32'h00402021; // 0040019c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h068: data = 32'h0c100257; // 004001a0: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h069: data = 32'h00000000; // 004001a4: SLL, REG[0]<=REG[0]<<0;
      10'h06a: data = 32'h2402000a; // 004001a8: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h06b: data = 32'hafc20024; // 004001ac: SW, RAM[REG[30]+36]<=REG[2];
      10'h06c: data = 32'hafc00028; // 004001b0: SW, RAM[REG[30]+40]<=REG[0];
      10'h06d: data = 32'h27c20024; // 004001b4: ADDIU, REG[2]<=REG[30]+36(=0x00000024);
      10'h06e: data = 32'h00402021; // 004001b8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h06f: data = 32'h0c100257; // 004001bc: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h070: data = 32'h00000000; // 004001c0: SLL, REG[0]<=REG[0]<<0;
      10'h071: data = 32'h27c20064; // 004001c4: ADDIU, REG[2]<=REG[30]+100(=0x00000064);
      10'h072: data = 32'h00402021; // 004001c8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h073: data = 32'h0c1000b8; // 004001cc: JAL, PC<=0x001000b8*4(=0x004002e0); REG[31]<=PC+4
      10'h074: data = 32'h00000000; // 004001d0: SLL, REG[0]<=REG[0]<<0;
      10'h075: data = 32'hafc20018; // 004001d4: SW, RAM[REG[30]+24]<=REG[2];
      10'h076: data = 32'h24020002; // 004001d8: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h077: data = 32'hafc2001c; // 004001dc: SW, RAM[REG[30]+28]<=REG[2];
      10'h078: data = 32'h081000a0; // 004001e0: J, PC<=0x001000a0*4(=0x00400280);
      10'h079: data = 32'h00000000; // 004001e4: SLL, REG[0]<=REG[0]<<0;
      10'h07a: data = 32'h8fc2001c; // 004001e8: LW, REG[2]<=RAM[REG[30]+28];
      10'h07b: data = 32'h8fc30020; // 004001ec: LW, REG[3]<=RAM[REG[30]+32];
      10'h07c: data = 32'h00021080; // 004001f0: SLL, REG[2]<=REG[2]<<2;
      10'h07d: data = 32'h00431021; // 004001f4: ADDU, REG[2]<=REG[2]+REG[3];
      10'h07e: data = 32'h8c430000; // 004001f8: LW, REG[3]<=RAM[REG[2]+0];
      10'h07f: data = 32'h24020001; // 004001fc: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h080: data = 32'h1462001b; // 00400200: BNE, PC<=(REG[3] != REG[2])?PC+4+27*4:PC+4;
      10'h081: data = 32'h00000000; // 00400204: SLL, REG[0]<=REG[0]<<0;
      10'h082: data = 32'h8fc2001c; // 00400208: LW, REG[2]<=RAM[REG[30]+28];
      10'h083: data = 32'h8fc3001c; // 0040020c: LW, REG[3]<=RAM[REG[30]+28];
      10'h084: data = 32'h00000000; // 00400210: SLL, REG[0]<=REG[0]<<0;
      10'h085: data = 32'h00431021; // 00400214: ADDU, REG[2]<=REG[2]+REG[3];
      10'h086: data = 32'hafc20014; // 00400218: SW, RAM[REG[30]+20]<=REG[2];
      10'h087: data = 32'h08100093; // 0040021c: J, PC<=0x00100093*4(=0x0040024c);
      10'h088: data = 32'h00000000; // 00400220: SLL, REG[0]<=REG[0]<<0;
      10'h089: data = 32'h8fc20014; // 00400224: LW, REG[2]<=RAM[REG[30]+20];
      10'h08a: data = 32'h8fc30020; // 00400228: LW, REG[3]<=RAM[REG[30]+32];
      10'h08b: data = 32'h00021080; // 0040022c: SLL, REG[2]<=REG[2]<<2;
      10'h08c: data = 32'h00431021; // 00400230: ADDU, REG[2]<=REG[2]+REG[3];
      10'h08d: data = 32'hac400000; // 00400234: SW, RAM[REG[2]+0]<=REG[0];
      10'h08e: data = 32'h8fc30014; // 00400238: LW, REG[3]<=RAM[REG[30]+20];
      10'h08f: data = 32'h8fc2001c; // 0040023c: LW, REG[2]<=RAM[REG[30]+28];
      10'h090: data = 32'h00000000; // 00400240: SLL, REG[0]<=REG[0]<<0;
      10'h091: data = 32'h00621021; // 00400244: ADDU, REG[2]<=REG[3]+REG[2];
      10'h092: data = 32'hafc20014; // 00400248: SW, RAM[REG[30]+20]<=REG[2];
      10'h093: data = 32'h8fc20014; // 0040024c: LW, REG[2]<=RAM[REG[30]+20];
      10'h094: data = 32'h8fc30018; // 00400250: LW, REG[3]<=RAM[REG[30]+24];
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h0062102b; // 00400258: SLTU, REG[2]<=(REG[3]<REG[2])?1:0;
      10'h097: data = 32'h1040fff1; // 0040025c: BEQ, PC<=(REG[2] == REG[0])?PC+4+65521*4:PC+4;
      10'h098: data = 32'h00000000; // 00400260: SLL, REG[0]<=REG[0]<<0;
      10'h099: data = 32'h8fc4001c; // 00400264: LW, REG[4]<=RAM[REG[30]+28];
      10'h09a: data = 32'h0c10014b; // 00400268: JAL, PC<=0x0010014b*4(=0x0040052c); REG[31]<=PC+4
      10'h09b: data = 32'h00000000; // 0040026c: SLL, REG[0]<=REG[0]<<0;
      10'h09c: data = 32'h8fc2001c; // 00400270: LW, REG[2]<=RAM[REG[30]+28];
      10'h09d: data = 32'h00000000; // 00400274: SLL, REG[0]<=REG[0]<<0;
      10'h09e: data = 32'h24420001; // 00400278: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h09f: data = 32'hafc2001c; // 0040027c: SW, RAM[REG[30]+28]<=REG[2];
      10'h0a0: data = 32'h8fc2001c; // 00400280: LW, REG[2]<=RAM[REG[30]+28];
      10'h0a1: data = 32'h8fc30018; // 00400284: LW, REG[3]<=RAM[REG[30]+24];
      10'h0a2: data = 32'h00000000; // 00400288: SLL, REG[0]<=REG[0]<<0;
      10'h0a3: data = 32'h0062102b; // 0040028c: SLTU, REG[2]<=(REG[3]<REG[2])?1:0;
      10'h0a4: data = 32'h1040ffd5; // 00400290: BEQ, PC<=(REG[2] == REG[0])?PC+4+65493*4:PC+4;
      10'h0a5: data = 32'h00000000; // 00400294: SLL, REG[0]<=REG[0]<<0;
      10'h0a6: data = 32'h2402000a; // 00400298: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h0a7: data = 32'hafc20024; // 0040029c: SW, RAM[REG[30]+36]<=REG[2];
      10'h0a8: data = 32'hafc00028; // 004002a0: SW, RAM[REG[30]+40]<=REG[0];
      10'h0a9: data = 32'h27c20024; // 004002a4: ADDIU, REG[2]<=REG[30]+36(=0x00000024);
      10'h0aa: data = 32'h00402021; // 004002a8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h0ab: data = 32'h0c100257; // 004002ac: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h0ac: data = 32'h00000000; // 004002b0: SLL, REG[0]<=REG[0]<<0;
      10'h0ad: data = 32'h08100046; // 004002b4: J, PC<=0x00100046*4(=0x00400118);
      10'h0ae: data = 32'h00000000; // 004002b8: SLL, REG[0]<=REG[0]<<0;
      10'h0af: data = 32'h27bdfff0; // 004002bc: ADDIU, REG[29]<=REG[29]+65520(=0x0000fff0);
      10'h0b0: data = 32'hafbe0008; // 004002c0: SW, RAM[REG[29]+8]<=REG[30];
      10'h0b1: data = 32'h03a0f021; // 004002c4: ADDU, REG[30]<=REG[29]+REG[0];
      10'h0b2: data = 32'hafc40010; // 004002c8: SW, RAM[REG[30]+16]<=REG[4];
      10'h0b3: data = 32'h03c0e821; // 004002cc: ADDU, REG[29]<=REG[30]+REG[0];
      10'h0b4: data = 32'h8fbe0008; // 004002d0: LW, REG[30]<=RAM[REG[29]+8];
      10'h0b5: data = 32'h27bd0010; // 004002d4: ADDIU, REG[29]<=REG[29]+16(=0x00000010);
      10'h0b6: data = 32'h03e00008; // 004002d8: JR, PC<=REG[31];
      10'h0b7: data = 32'h00000000; // 004002dc: SLL, REG[0]<=REG[0]<<0;
      10'h0b8: data = 32'h27bdffe8; // 004002e0: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h0b9: data = 32'hafbe0010; // 004002e4: SW, RAM[REG[29]+16]<=REG[30];
      10'h0ba: data = 32'h03a0f021; // 004002e8: ADDU, REG[30]<=REG[29]+REG[0];
      10'h0bb: data = 32'hafc40018; // 004002ec: SW, RAM[REG[30]+24]<=REG[4];
      10'h0bc: data = 32'h8fc20018; // 004002f0: LW, REG[2]<=RAM[REG[30]+24];
      10'h0bd: data = 32'h00000000; // 004002f4: SLL, REG[0]<=REG[0]<<0;
      10'h0be: data = 32'hafc20008; // 004002f8: SW, RAM[REG[30]+8]<=REG[2];
      10'h0bf: data = 32'hafc00004; // 004002fc: SW, RAM[REG[30]+4]<=REG[0];
      10'h0c0: data = 32'h081000ca; // 00400300: J, PC<=0x001000ca*4(=0x00400328);
      10'h0c1: data = 32'h00000000; // 00400304: SLL, REG[0]<=REG[0]<<0;
      10'h0c2: data = 32'h8fc20008; // 00400308: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c3: data = 32'h00000000; // 0040030c: SLL, REG[0]<=REG[0]<<0;
      10'h0c4: data = 32'h24420004; // 00400310: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h0c5: data = 32'hafc20008; // 00400314: SW, RAM[REG[30]+8]<=REG[2];
      10'h0c6: data = 32'h8fc20004; // 00400318: LW, REG[2]<=RAM[REG[30]+4];
      10'h0c7: data = 32'h00000000; // 0040031c: SLL, REG[0]<=REG[0]<<0;
      10'h0c8: data = 32'h24420001; // 00400320: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h0c9: data = 32'hafc20004; // 00400324: SW, RAM[REG[30]+4]<=REG[2];
      10'h0ca: data = 32'h8fc20008; // 00400328: LW, REG[2]<=RAM[REG[30]+8];
      10'h0cb: data = 32'h00000000; // 0040032c: SLL, REG[0]<=REG[0]<<0;
      10'h0cc: data = 32'h8c420000; // 00400330: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cd: data = 32'h00000000; // 00400334: SLL, REG[0]<=REG[0]<<0;
      10'h0ce: data = 32'h1440fff3; // 00400338: BNE, PC<=(REG[2] != REG[0])?PC+4+65523*4:PC+4;
      10'h0cf: data = 32'h00000000; // 0040033c: SLL, REG[0]<=REG[0]<<0;
      10'h0d0: data = 32'hafc00000; // 00400340: SW, RAM[REG[30]+0]<=REG[0];
      10'h0d1: data = 32'h8fc20018; // 00400344: LW, REG[2]<=RAM[REG[30]+24];
      10'h0d2: data = 32'h00000000; // 00400348: SLL, REG[0]<=REG[0]<<0;
      10'h0d3: data = 32'hafc20008; // 0040034c: SW, RAM[REG[30]+8]<=REG[2];
      10'h0d4: data = 32'h8fc30004; // 00400350: LW, REG[3]<=RAM[REG[30]+4];
      10'h0d5: data = 32'h24020001; // 00400354: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0d6: data = 32'h14620009; // 00400358: BNE, PC<=(REG[3] != REG[2])?PC+4+9*4:PC+4;
      10'h0d7: data = 32'h00000000; // 0040035c: SLL, REG[0]<=REG[0]<<0;
      10'h0d8: data = 32'h8fc20008; // 00400360: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d9: data = 32'h00000000; // 00400364: SLL, REG[0]<=REG[0]<<0;
      10'h0da: data = 32'h8c420000; // 00400368: LW, REG[2]<=RAM[REG[2]+0];
      10'h0db: data = 32'h00000000; // 0040036c: SLL, REG[0]<=REG[0]<<0;
      10'h0dc: data = 32'h2442ffd0; // 00400370: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h0dd: data = 32'hafc20000; // 00400374: SW, RAM[REG[30]+0]<=REG[2];
      10'h0de: data = 32'h08100145; // 00400378: J, PC<=0x00100145*4(=0x00400514);
      10'h0df: data = 32'h00000000; // 0040037c: SLL, REG[0]<=REG[0]<<0;
      10'h0e0: data = 32'h8fc30004; // 00400380: LW, REG[3]<=RAM[REG[30]+4];
      10'h0e1: data = 32'h24020002; // 00400384: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h0e2: data = 32'h14620024; // 00400388: BNE, PC<=(REG[3] != REG[2])?PC+4+36*4:PC+4;
      10'h0e3: data = 32'h00000000; // 0040038c: SLL, REG[0]<=REG[0]<<0;
      10'h0e4: data = 32'hafc00004; // 00400390: SW, RAM[REG[30]+4]<=REG[0];
      10'h0e5: data = 32'h081000ef; // 00400394: J, PC<=0x001000ef*4(=0x004003bc);
      10'h0e6: data = 32'h00000000; // 00400398: SLL, REG[0]<=REG[0]<<0;
      10'h0e7: data = 32'h8fc20000; // 0040039c: LW, REG[2]<=RAM[REG[30]+0];
      10'h0e8: data = 32'h00000000; // 004003a0: SLL, REG[0]<=REG[0]<<0;
      10'h0e9: data = 32'h2442000a; // 004003a4: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h0ea: data = 32'hafc20000; // 004003a8: SW, RAM[REG[30]+0]<=REG[2];
      10'h0eb: data = 32'h8fc20004; // 004003ac: LW, REG[2]<=RAM[REG[30]+4];
      10'h0ec: data = 32'h00000000; // 004003b0: SLL, REG[0]<=REG[0]<<0;
      10'h0ed: data = 32'h24420001; // 004003b4: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h0ee: data = 32'hafc20004; // 004003b8: SW, RAM[REG[30]+4]<=REG[2];
      10'h0ef: data = 32'h8fc20008; // 004003bc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f0: data = 32'h00000000; // 004003c0: SLL, REG[0]<=REG[0]<<0;
      10'h0f1: data = 32'h8c420000; // 004003c4: LW, REG[2]<=RAM[REG[2]+0];
      10'h0f2: data = 32'h00000000; // 004003c8: SLL, REG[0]<=REG[0]<<0;
      10'h0f3: data = 32'h2443ffd0; // 004003cc: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h0f4: data = 32'h8fc20004; // 004003d0: LW, REG[2]<=RAM[REG[30]+4];
      10'h0f5: data = 32'h00000000; // 004003d4: SLL, REG[0]<=REG[0]<<0;
      10'h0f6: data = 32'h0043102b; // 004003d8: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h0f7: data = 32'h1440ffef; // 004003dc: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h0f8: data = 32'h00000000; // 004003e0: SLL, REG[0]<=REG[0]<<0;
      10'h0f9: data = 32'h8fc20008; // 004003e4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0fa: data = 32'h00000000; // 004003e8: SLL, REG[0]<=REG[0]<<0;
      10'h0fb: data = 32'h24420004; // 004003ec: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h0fc: data = 32'hafc20008; // 004003f0: SW, RAM[REG[30]+8]<=REG[2];
      10'h0fd: data = 32'h8fc20008; // 004003f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0fe: data = 32'h00000000; // 004003f8: SLL, REG[0]<=REG[0]<<0;
      10'h0ff: data = 32'h8c430000; // 004003fc: LW, REG[3]<=RAM[REG[2]+0];
      10'h100: data = 32'h8fc20000; // 00400400: LW, REG[2]<=RAM[REG[30]+0];
      10'h101: data = 32'h00000000; // 00400404: SLL, REG[0]<=REG[0]<<0;
      10'h102: data = 32'h00621021; // 00400408: ADDU, REG[2]<=REG[3]+REG[2];
      10'h103: data = 32'h2442ffd0; // 0040040c: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h104: data = 32'hafc20000; // 00400410: SW, RAM[REG[30]+0]<=REG[2];
      10'h105: data = 32'h08100145; // 00400414: J, PC<=0x00100145*4(=0x00400514);
      10'h106: data = 32'h00000000; // 00400418: SLL, REG[0]<=REG[0]<<0;
      10'h107: data = 32'h8fc30004; // 0040041c: LW, REG[3]<=RAM[REG[30]+4];
      10'h108: data = 32'h24020003; // 00400420: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h109: data = 32'h1462003b; // 00400424: BNE, PC<=(REG[3] != REG[2])?PC+4+59*4:PC+4;
      10'h10a: data = 32'h00000000; // 00400428: SLL, REG[0]<=REG[0]<<0;
      10'h10b: data = 32'hafc00004; // 0040042c: SW, RAM[REG[30]+4]<=REG[0];
      10'h10c: data = 32'h08100116; // 00400430: J, PC<=0x00100116*4(=0x00400458);
      10'h10d: data = 32'h00000000; // 00400434: SLL, REG[0]<=REG[0]<<0;
      10'h10e: data = 32'h8fc20000; // 00400438: LW, REG[2]<=RAM[REG[30]+0];
      10'h10f: data = 32'h00000000; // 0040043c: SLL, REG[0]<=REG[0]<<0;
      10'h110: data = 32'h24420064; // 00400440: ADDIU, REG[2]<=REG[2]+100(=0x00000064);
      10'h111: data = 32'hafc20000; // 00400444: SW, RAM[REG[30]+0]<=REG[2];
      10'h112: data = 32'h8fc20004; // 00400448: LW, REG[2]<=RAM[REG[30]+4];
      10'h113: data = 32'h00000000; // 0040044c: SLL, REG[0]<=REG[0]<<0;
      10'h114: data = 32'h24420001; // 00400450: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h115: data = 32'hafc20004; // 00400454: SW, RAM[REG[30]+4]<=REG[2];
      10'h116: data = 32'h8fc20008; // 00400458: LW, REG[2]<=RAM[REG[30]+8];
      10'h117: data = 32'h00000000; // 0040045c: SLL, REG[0]<=REG[0]<<0;
      10'h118: data = 32'h8c420000; // 00400460: LW, REG[2]<=RAM[REG[2]+0];
      10'h119: data = 32'h00000000; // 00400464: SLL, REG[0]<=REG[0]<<0;
      10'h11a: data = 32'h2443ffd0; // 00400468: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h11b: data = 32'h8fc20004; // 0040046c: LW, REG[2]<=RAM[REG[30]+4];
      10'h11c: data = 32'h00000000; // 00400470: SLL, REG[0]<=REG[0]<<0;
      10'h11d: data = 32'h0043102b; // 00400474: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h11e: data = 32'h1440ffef; // 00400478: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h11f: data = 32'h00000000; // 0040047c: SLL, REG[0]<=REG[0]<<0;
      10'h120: data = 32'h8fc20008; // 00400480: LW, REG[2]<=RAM[REG[30]+8];
      10'h121: data = 32'h00000000; // 00400484: SLL, REG[0]<=REG[0]<<0;
      10'h122: data = 32'h24420004; // 00400488: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h123: data = 32'hafc20008; // 0040048c: SW, RAM[REG[30]+8]<=REG[2];
      10'h124: data = 32'hafc00004; // 00400490: SW, RAM[REG[30]+4]<=REG[0];
      10'h125: data = 32'h0810012f; // 00400494: J, PC<=0x0010012f*4(=0x004004bc);
      10'h126: data = 32'h00000000; // 00400498: SLL, REG[0]<=REG[0]<<0;
      10'h127: data = 32'h8fc20000; // 0040049c: LW, REG[2]<=RAM[REG[30]+0];
      10'h128: data = 32'h00000000; // 004004a0: SLL, REG[0]<=REG[0]<<0;
      10'h129: data = 32'h2442000a; // 004004a4: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h12a: data = 32'hafc20000; // 004004a8: SW, RAM[REG[30]+0]<=REG[2];
      10'h12b: data = 32'h8fc20004; // 004004ac: LW, REG[2]<=RAM[REG[30]+4];
      10'h12c: data = 32'h00000000; // 004004b0: SLL, REG[0]<=REG[0]<<0;
      10'h12d: data = 32'h24420001; // 004004b4: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h12e: data = 32'hafc20004; // 004004b8: SW, RAM[REG[30]+4]<=REG[2];
      10'h12f: data = 32'h8fc20008; // 004004bc: LW, REG[2]<=RAM[REG[30]+8];
      10'h130: data = 32'h00000000; // 004004c0: SLL, REG[0]<=REG[0]<<0;
      10'h131: data = 32'h8c420000; // 004004c4: LW, REG[2]<=RAM[REG[2]+0];
      10'h132: data = 32'h00000000; // 004004c8: SLL, REG[0]<=REG[0]<<0;
      10'h133: data = 32'h2443ffd0; // 004004cc: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h134: data = 32'h8fc20004; // 004004d0: LW, REG[2]<=RAM[REG[30]+4];
      10'h135: data = 32'h00000000; // 004004d4: SLL, REG[0]<=REG[0]<<0;
      10'h136: data = 32'h0043102b; // 004004d8: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h137: data = 32'h1440ffef; // 004004dc: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h138: data = 32'h00000000; // 004004e0: SLL, REG[0]<=REG[0]<<0;
      10'h139: data = 32'h8fc20008; // 004004e4: LW, REG[2]<=RAM[REG[30]+8];
      10'h13a: data = 32'h00000000; // 004004e8: SLL, REG[0]<=REG[0]<<0;
      10'h13b: data = 32'h24420004; // 004004ec: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h13c: data = 32'hafc20008; // 004004f0: SW, RAM[REG[30]+8]<=REG[2];
      10'h13d: data = 32'h8fc20008; // 004004f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h13e: data = 32'h00000000; // 004004f8: SLL, REG[0]<=REG[0]<<0;
      10'h13f: data = 32'h8c430000; // 004004fc: LW, REG[3]<=RAM[REG[2]+0];
      10'h140: data = 32'h8fc20000; // 00400500: LW, REG[2]<=RAM[REG[30]+0];
      10'h141: data = 32'h00000000; // 00400504: SLL, REG[0]<=REG[0]<<0;
      10'h142: data = 32'h00621021; // 00400508: ADDU, REG[2]<=REG[3]+REG[2];
      10'h143: data = 32'h2442ffd0; // 0040050c: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h144: data = 32'hafc20000; // 00400510: SW, RAM[REG[30]+0]<=REG[2];
      10'h145: data = 32'h8fc20000; // 00400514: LW, REG[2]<=RAM[REG[30]+0];
      10'h146: data = 32'h03c0e821; // 00400518: ADDU, REG[29]<=REG[30]+REG[0];
      10'h147: data = 32'h8fbe0010; // 0040051c: LW, REG[30]<=RAM[REG[29]+16];
      10'h148: data = 32'h27bd0018; // 00400520: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h149: data = 32'h03e00008; // 00400524: JR, PC<=REG[31];
      10'h14a: data = 32'h00000000; // 00400528: SLL, REG[0]<=REG[0]<<0;
      10'h14b: data = 32'h27bdffd0; // 0040052c: ADDIU, REG[29]<=REG[29]+65488(=0x0000ffd0);
      10'h14c: data = 32'hafbf002c; // 00400530: SW, RAM[REG[29]+44]<=REG[31];
      10'h14d: data = 32'hafbe0028; // 00400534: SW, RAM[REG[29]+40]<=REG[30];
      10'h14e: data = 32'h03a0f021; // 00400538: ADDU, REG[30]<=REG[29]+REG[0];
      10'h14f: data = 32'hafc40030; // 0040053c: SW, RAM[REG[30]+48]<=REG[4];
      10'h150: data = 32'hafc00010; // 00400540: SW, RAM[REG[30]+16]<=REG[0];
      10'h151: data = 32'h0810015b; // 00400544: J, PC<=0x0010015b*4(=0x0040056c);
      10'h152: data = 32'h00000000; // 00400548: SLL, REG[0]<=REG[0]<<0;
      10'h153: data = 32'h8fc20030; // 0040054c: LW, REG[2]<=RAM[REG[30]+48];
      10'h154: data = 32'h00000000; // 00400550: SLL, REG[0]<=REG[0]<<0;
      10'h155: data = 32'h2442fff6; // 00400554: ADDIU, REG[2]<=REG[2]+65526(=0x0000fff6);
      10'h156: data = 32'hafc20030; // 00400558: SW, RAM[REG[30]+48]<=REG[2];
      10'h157: data = 32'h8fc20010; // 0040055c: LW, REG[2]<=RAM[REG[30]+16];
      10'h158: data = 32'h00000000; // 00400560: SLL, REG[0]<=REG[0]<<0;
      10'h159: data = 32'h24420001; // 00400564: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h15a: data = 32'hafc20010; // 00400568: SW, RAM[REG[30]+16]<=REG[2];
      10'h15b: data = 32'h8fc20030; // 0040056c: LW, REG[2]<=RAM[REG[30]+48];
      10'h15c: data = 32'h00000000; // 00400570: SLL, REG[0]<=REG[0]<<0;
      10'h15d: data = 32'h2c42000a; // 00400574: SLTIU, REG[2]<=(REG[2]<10(=0x0000000a))?1:0;
      10'h15e: data = 32'h1040fff4; // 00400578: BEQ, PC<=(REG[2] == REG[0])?PC+4+65524*4:PC+4;
      10'h15f: data = 32'h00000000; // 0040057c: SLL, REG[0]<=REG[0]<<0;
      10'h160: data = 32'h8fc20010; // 00400580: LW, REG[2]<=RAM[REG[30]+16];
      10'h161: data = 32'h00000000; // 00400584: SLL, REG[0]<=REG[0]<<0;
      10'h162: data = 32'h24420030; // 00400588: ADDIU, REG[2]<=REG[2]+48(=0x00000030);
      10'h163: data = 32'hafc20014; // 0040058c: SW, RAM[REG[30]+20]<=REG[2];
      10'h164: data = 32'h8fc20030; // 00400590: LW, REG[2]<=RAM[REG[30]+48];
      10'h165: data = 32'h00000000; // 00400594: SLL, REG[0]<=REG[0]<<0;
      10'h166: data = 32'h24420030; // 00400598: ADDIU, REG[2]<=REG[2]+48(=0x00000030);
      10'h167: data = 32'hafc20018; // 0040059c: SW, RAM[REG[30]+24]<=REG[2];
      10'h168: data = 32'h24020020; // 004005a0: ADDIU, REG[2]<=REG[0]+32(=0x00000020);
      10'h169: data = 32'hafc2001c; // 004005a4: SW, RAM[REG[30]+28]<=REG[2];
      10'h16a: data = 32'hafc00020; // 004005a8: SW, RAM[REG[30]+32]<=REG[0];
      10'h16b: data = 32'h27c20014; // 004005ac: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h16c: data = 32'h00402021; // 004005b0: ADDU, REG[4]<=REG[2]+REG[0];
      10'h16d: data = 32'h0c100257; // 004005b4: JAL, PC<=0x00100257*4(=0x0040095c); REG[31]<=PC+4
      10'h16e: data = 32'h00000000; // 004005b8: SLL, REG[0]<=REG[0]<<0;
      10'h16f: data = 32'h03c0e821; // 004005bc: ADDU, REG[29]<=REG[30]+REG[0];
      10'h170: data = 32'h8fbf002c; // 004005c0: LW, REG[31]<=RAM[REG[29]+44];
      10'h171: data = 32'h8fbe0028; // 004005c4: LW, REG[30]<=RAM[REG[29]+40];
      10'h172: data = 32'h27bd0030; // 004005c8: ADDIU, REG[29]<=REG[29]+48(=0x00000030);
      10'h173: data = 32'h03e00008; // 004005cc: JR, PC<=REG[31];
      10'h174: data = 32'h00000000; // 004005d0: SLL, REG[0]<=REG[0]<<0;
      10'h175: data = 32'h27bdfff8; // 004005d4: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h176: data = 32'hafbe0000; // 004005d8: SW, RAM[REG[29]+0]<=REG[30];
      10'h177: data = 32'h03a0f021; // 004005dc: ADDU, REG[30]<=REG[29]+REG[0];
      10'h178: data = 32'hafc40008; // 004005e0: SW, RAM[REG[30]+8]<=REG[4];
      10'h179: data = 32'h24020308; // 004005e4: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h17a: data = 32'hac400000; // 004005e8: SW, RAM[REG[2]+0]<=REG[0];
      10'h17b: data = 32'h2403030c; // 004005ec: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h17c: data = 32'h24020001; // 004005f0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h17d: data = 32'hac620000; // 004005f4: SW, RAM[REG[3]+0]<=REG[2];
      10'h17e: data = 32'h24030308; // 004005f8: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h17f: data = 32'h24020001; // 004005fc: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h180: data = 32'hac620000; // 00400600: SW, RAM[REG[3]+0]<=REG[2];
      10'h181: data = 32'h24020308; // 00400604: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h182: data = 32'hac400000; // 00400608: SW, RAM[REG[2]+0]<=REG[0];
      10'h183: data = 32'h24030308; // 0040060c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h184: data = 32'h24020001; // 00400610: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h185: data = 32'hac620000; // 00400614: SW, RAM[REG[3]+0]<=REG[2];
      10'h186: data = 32'h0810018d; // 00400618: J, PC<=0x0010018d*4(=0x00400634);
      10'h187: data = 32'h00000000; // 0040061c: SLL, REG[0]<=REG[0]<<0;
      10'h188: data = 32'h24020308; // 00400620: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h189: data = 32'hac400000; // 00400624: SW, RAM[REG[2]+0]<=REG[0];
      10'h18a: data = 32'h24030308; // 00400628: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h18b: data = 32'h24020001; // 0040062c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h18c: data = 32'hac620000; // 00400630: SW, RAM[REG[3]+0]<=REG[2];
      10'h18d: data = 32'h24020310; // 00400634: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h18e: data = 32'h8c430000; // 00400638: LW, REG[3]<=RAM[REG[2]+0];
      10'h18f: data = 32'h2402ffff; // 0040063c: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h190: data = 32'h1062fff7; // 00400640: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h191: data = 32'h00000000; // 00400644: SLL, REG[0]<=REG[0]<<0;
      10'h192: data = 32'h0810023b; // 00400648: J, PC<=0x0010023b*4(=0x004008ec);
      10'h193: data = 32'h00000000; // 0040064c: SLL, REG[0]<=REG[0]<<0;
      10'h194: data = 32'h8fc20008; // 00400650: LW, REG[2]<=RAM[REG[30]+8];
      10'h195: data = 32'h00000000; // 00400654: SLL, REG[0]<=REG[0]<<0;
      10'h196: data = 32'h8c420000; // 00400658: LW, REG[2]<=RAM[REG[2]+0];
      10'h197: data = 32'h00000000; // 0040065c: SLL, REG[0]<=REG[0]<<0;
      10'h198: data = 32'h10400012; // 00400660: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h199: data = 32'h00000000; // 00400664: SLL, REG[0]<=REG[0]<<0;
      10'h19a: data = 32'h8fc20008; // 00400668: LW, REG[2]<=RAM[REG[30]+8];
      10'h19b: data = 32'h00000000; // 0040066c: SLL, REG[0]<=REG[0]<<0;
      10'h19c: data = 32'h8c420000; // 00400670: LW, REG[2]<=RAM[REG[2]+0];
      10'h19d: data = 32'h00000000; // 00400674: SLL, REG[0]<=REG[0]<<0;
      10'h19e: data = 32'h2c42001b; // 00400678: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h19f: data = 32'h1040000b; // 0040067c: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h1a0: data = 32'h00000000; // 00400680: SLL, REG[0]<=REG[0]<<0;
      10'h1a1: data = 32'h8fc20008; // 00400684: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a2: data = 32'h00000000; // 00400688: SLL, REG[0]<=REG[0]<<0;
      10'h1a3: data = 32'h8c420000; // 0040068c: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a4: data = 32'h00000000; // 00400690: SLL, REG[0]<=REG[0]<<0;
      10'h1a5: data = 32'h24430040; // 00400694: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h1a6: data = 32'h8fc20008; // 00400698: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a7: data = 32'h00000000; // 0040069c: SLL, REG[0]<=REG[0]<<0;
      10'h1a8: data = 32'hac430000; // 004006a0: SW, RAM[REG[2]+0]<=REG[3];
      10'h1a9: data = 32'h08100232; // 004006a4: J, PC<=0x00100232*4(=0x004008c8);
      10'h1aa: data = 32'h00000000; // 004006a8: SLL, REG[0]<=REG[0]<<0;
      10'h1ab: data = 32'h8fc20008; // 004006ac: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ac: data = 32'h00000000; // 004006b0: SLL, REG[0]<=REG[0]<<0;
      10'h1ad: data = 32'h8c420000; // 004006b4: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ae: data = 32'h00000000; // 004006b8: SLL, REG[0]<=REG[0]<<0;
      10'h1af: data = 32'h2c420030; // 004006bc: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1b0: data = 32'h14400010; // 004006c0: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1b1: data = 32'h00000000; // 004006c4: SLL, REG[0]<=REG[0]<<0;
      10'h1b2: data = 32'h8fc20008; // 004006c8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b3: data = 32'h00000000; // 004006cc: SLL, REG[0]<=REG[0]<<0;
      10'h1b4: data = 32'h8c420000; // 004006d0: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b5: data = 32'h00000000; // 004006d4: SLL, REG[0]<=REG[0]<<0;
      10'h1b6: data = 32'h2c42003a; // 004006d8: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h1b7: data = 32'h10400009; // 004006dc: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1b8: data = 32'h00000000; // 004006e0: SLL, REG[0]<=REG[0]<<0;
      10'h1b9: data = 32'h8fc20008; // 004006e4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ba: data = 32'h00000000; // 004006e8: SLL, REG[0]<=REG[0]<<0;
      10'h1bb: data = 32'h8c430000; // 004006ec: LW, REG[3]<=RAM[REG[2]+0];
      10'h1bc: data = 32'h8fc20008; // 004006f0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1bd: data = 32'h00000000; // 004006f4: SLL, REG[0]<=REG[0]<<0;
      10'h1be: data = 32'hac430000; // 004006f8: SW, RAM[REG[2]+0]<=REG[3];
      10'h1bf: data = 32'h08100232; // 004006fc: J, PC<=0x00100232*4(=0x004008c8);
      10'h1c0: data = 32'h00000000; // 00400700: SLL, REG[0]<=REG[0]<<0;
      10'h1c1: data = 32'h8fc20008; // 00400704: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c2: data = 32'h00000000; // 00400708: SLL, REG[0]<=REG[0]<<0;
      10'h1c3: data = 32'h8c420000; // 0040070c: LW, REG[2]<=RAM[REG[2]+0];
      10'h1c4: data = 32'h00000000; // 00400710: SLL, REG[0]<=REG[0]<<0;
      10'h1c5: data = 32'h14400006; // 00400714: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h1c6: data = 32'h00000000; // 00400718: SLL, REG[0]<=REG[0]<<0;
      10'h1c7: data = 32'h8fc30008; // 0040071c: LW, REG[3]<=RAM[REG[30]+8];
      10'h1c8: data = 32'h24020040; // 00400720: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h1c9: data = 32'hac620000; // 00400724: SW, RAM[REG[3]+0]<=REG[2];
      10'h1ca: data = 32'h08100232; // 00400728: J, PC<=0x00100232*4(=0x004008c8);
      10'h1cb: data = 32'h00000000; // 0040072c: SLL, REG[0]<=REG[0]<<0;
      10'h1cc: data = 32'h8fc20008; // 00400730: LW, REG[2]<=RAM[REG[30]+8];
      10'h1cd: data = 32'h00000000; // 00400734: SLL, REG[0]<=REG[0]<<0;
      10'h1ce: data = 32'h8c430000; // 00400738: LW, REG[3]<=RAM[REG[2]+0];
      10'h1cf: data = 32'h2402001b; // 0040073c: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h1d0: data = 32'h14620006; // 00400740: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1d1: data = 32'h00000000; // 00400744: SLL, REG[0]<=REG[0]<<0;
      10'h1d2: data = 32'h8fc30008; // 00400748: LW, REG[3]<=RAM[REG[30]+8];
      10'h1d3: data = 32'h2402005b; // 0040074c: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h1d4: data = 32'hac620000; // 00400750: SW, RAM[REG[3]+0]<=REG[2];
      10'h1d5: data = 32'h08100232; // 00400754: J, PC<=0x00100232*4(=0x004008c8);
      10'h1d6: data = 32'h00000000; // 00400758: SLL, REG[0]<=REG[0]<<0;
      10'h1d7: data = 32'h8fc20008; // 0040075c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1d8: data = 32'h00000000; // 00400760: SLL, REG[0]<=REG[0]<<0;
      10'h1d9: data = 32'h8c430000; // 00400764: LW, REG[3]<=RAM[REG[2]+0];
      10'h1da: data = 32'h2402001d; // 00400768: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h1db: data = 32'h14620006; // 0040076c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1dc: data = 32'h00000000; // 00400770: SLL, REG[0]<=REG[0]<<0;
      10'h1dd: data = 32'h8fc30008; // 00400774: LW, REG[3]<=RAM[REG[30]+8];
      10'h1de: data = 32'h2402005d; // 00400778: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h1df: data = 32'hac620000; // 0040077c: SW, RAM[REG[3]+0]<=REG[2];
      10'h1e0: data = 32'h08100232; // 00400780: J, PC<=0x00100232*4(=0x004008c8);
      10'h1e1: data = 32'h00000000; // 00400784: SLL, REG[0]<=REG[0]<<0;
      10'h1e2: data = 32'h8fc20008; // 00400788: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e3: data = 32'h00000000; // 0040078c: SLL, REG[0]<=REG[0]<<0;
      10'h1e4: data = 32'h8c420000; // 00400790: LW, REG[2]<=RAM[REG[2]+0];
      10'h1e5: data = 32'h00000000; // 00400794: SLL, REG[0]<=REG[0]<<0;
      10'h1e6: data = 32'h2c420020; // 00400798: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h1e7: data = 32'h14400010; // 0040079c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1e8: data = 32'h00000000; // 004007a0: SLL, REG[0]<=REG[0]<<0;
      10'h1e9: data = 32'h8fc20008; // 004007a4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ea: data = 32'h00000000; // 004007a8: SLL, REG[0]<=REG[0]<<0;
      10'h1eb: data = 32'h8c420000; // 004007ac: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ec: data = 32'h00000000; // 004007b0: SLL, REG[0]<=REG[0]<<0;
      10'h1ed: data = 32'h2c420030; // 004007b4: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1ee: data = 32'h10400009; // 004007b8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1ef: data = 32'h00000000; // 004007bc: SLL, REG[0]<=REG[0]<<0;
      10'h1f0: data = 32'h8fc20008; // 004007c0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f1: data = 32'h00000000; // 004007c4: SLL, REG[0]<=REG[0]<<0;
      10'h1f2: data = 32'h8c430000; // 004007c8: LW, REG[3]<=RAM[REG[2]+0];
      10'h1f3: data = 32'h8fc20008; // 004007cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f4: data = 32'h00000000; // 004007d0: SLL, REG[0]<=REG[0]<<0;
      10'h1f5: data = 32'hac430000; // 004007d4: SW, RAM[REG[2]+0]<=REG[3];
      10'h1f6: data = 32'h08100232; // 004007d8: J, PC<=0x00100232*4(=0x004008c8);
      10'h1f7: data = 32'h00000000; // 004007dc: SLL, REG[0]<=REG[0]<<0;
      10'h1f8: data = 32'h8fc20008; // 004007e0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f9: data = 32'h00000000; // 004007e4: SLL, REG[0]<=REG[0]<<0;
      10'h1fa: data = 32'h8c430000; // 004007e8: LW, REG[3]<=RAM[REG[2]+0];
      10'h1fb: data = 32'h2402003a; // 004007ec: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h1fc: data = 32'h14620006; // 004007f0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1fd: data = 32'h00000000; // 004007f4: SLL, REG[0]<=REG[0]<<0;
      10'h1fe: data = 32'h8fc30008; // 004007f8: LW, REG[3]<=RAM[REG[30]+8];
      10'h1ff: data = 32'h2402003f; // 004007fc: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h200: data = 32'hac620000; // 00400800: SW, RAM[REG[3]+0]<=REG[2];
      10'h201: data = 32'h08100232; // 00400804: J, PC<=0x00100232*4(=0x004008c8);
      10'h202: data = 32'h00000000; // 00400808: SLL, REG[0]<=REG[0]<<0;
      10'h203: data = 32'h8fc20008; // 0040080c: LW, REG[2]<=RAM[REG[30]+8];
      10'h204: data = 32'h00000000; // 00400810: SLL, REG[0]<=REG[0]<<0;
      10'h205: data = 32'h8c430000; // 00400814: LW, REG[3]<=RAM[REG[2]+0];
      10'h206: data = 32'h2402003b; // 00400818: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h207: data = 32'h14620006; // 0040081c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h208: data = 32'h00000000; // 00400820: SLL, REG[0]<=REG[0]<<0;
      10'h209: data = 32'h8fc30008; // 00400824: LW, REG[3]<=RAM[REG[30]+8];
      10'h20a: data = 32'h2402003d; // 00400828: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h20b: data = 32'hac620000; // 0040082c: SW, RAM[REG[3]+0]<=REG[2];
      10'h20c: data = 32'h08100232; // 00400830: J, PC<=0x00100232*4(=0x004008c8);
      10'h20d: data = 32'h00000000; // 00400834: SLL, REG[0]<=REG[0]<<0;
      10'h20e: data = 32'h8fc20008; // 00400838: LW, REG[2]<=RAM[REG[30]+8];
      10'h20f: data = 32'h00000000; // 0040083c: SLL, REG[0]<=REG[0]<<0;
      10'h210: data = 32'h8c430000; // 00400840: LW, REG[3]<=RAM[REG[2]+0];
      10'h211: data = 32'h2402003c; // 00400844: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h212: data = 32'h14620006; // 00400848: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h213: data = 32'h00000000; // 0040084c: SLL, REG[0]<=REG[0]<<0;
      10'h214: data = 32'h8fc30008; // 00400850: LW, REG[3]<=RAM[REG[30]+8];
      10'h215: data = 32'h2402003b; // 00400854: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h216: data = 32'hac620000; // 00400858: SW, RAM[REG[3]+0]<=REG[2];
      10'h217: data = 32'h08100232; // 0040085c: J, PC<=0x00100232*4(=0x004008c8);
      10'h218: data = 32'h00000000; // 00400860: SLL, REG[0]<=REG[0]<<0;
      10'h219: data = 32'h8fc20008; // 00400864: LW, REG[2]<=RAM[REG[30]+8];
      10'h21a: data = 32'h00000000; // 00400868: SLL, REG[0]<=REG[0]<<0;
      10'h21b: data = 32'h8c430000; // 0040086c: LW, REG[3]<=RAM[REG[2]+0];
      10'h21c: data = 32'h2402003d; // 00400870: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h21d: data = 32'h14620006; // 00400874: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h21e: data = 32'h00000000; // 00400878: SLL, REG[0]<=REG[0]<<0;
      10'h21f: data = 32'h8fc30008; // 0040087c: LW, REG[3]<=RAM[REG[30]+8];
      10'h220: data = 32'h2402003a; // 00400880: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h221: data = 32'hac620000; // 00400884: SW, RAM[REG[3]+0]<=REG[2];
      10'h222: data = 32'h08100232; // 00400888: J, PC<=0x00100232*4(=0x004008c8);
      10'h223: data = 32'h00000000; // 0040088c: SLL, REG[0]<=REG[0]<<0;
      10'h224: data = 32'h8fc20008; // 00400890: LW, REG[2]<=RAM[REG[30]+8];
      10'h225: data = 32'h00000000; // 00400894: SLL, REG[0]<=REG[0]<<0;
      10'h226: data = 32'h8c430000; // 00400898: LW, REG[3]<=RAM[REG[2]+0];
      10'h227: data = 32'h2402003e; // 0040089c: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h228: data = 32'h14620006; // 004008a0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h229: data = 32'h00000000; // 004008a4: SLL, REG[0]<=REG[0]<<0;
      10'h22a: data = 32'h8fc30008; // 004008a8: LW, REG[3]<=RAM[REG[30]+8];
      10'h22b: data = 32'h2402000a; // 004008ac: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h22c: data = 32'hac620000; // 004008b0: SW, RAM[REG[3]+0]<=REG[2];
      10'h22d: data = 32'h08100232; // 004008b4: J, PC<=0x00100232*4(=0x004008c8);
      10'h22e: data = 32'h00000000; // 004008b8: SLL, REG[0]<=REG[0]<<0;
      10'h22f: data = 32'h8fc30008; // 004008bc: LW, REG[3]<=RAM[REG[30]+8];
      10'h230: data = 32'h24020040; // 004008c0: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h231: data = 32'hac620000; // 004008c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h232: data = 32'h24020308; // 004008c8: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h233: data = 32'hac400000; // 004008cc: SW, RAM[REG[2]+0]<=REG[0];
      10'h234: data = 32'h24030308; // 004008d0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h235: data = 32'h24020001; // 004008d4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h236: data = 32'hac620000; // 004008d8: SW, RAM[REG[3]+0]<=REG[2];
      10'h237: data = 32'h8fc20008; // 004008dc: LW, REG[2]<=RAM[REG[30]+8];
      10'h238: data = 32'h00000000; // 004008e0: SLL, REG[0]<=REG[0]<<0;
      10'h239: data = 32'h24420004; // 004008e4: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h23a: data = 32'hafc20008; // 004008e8: SW, RAM[REG[30]+8]<=REG[2];
      10'h23b: data = 32'h24020310; // 004008ec: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h23c: data = 32'h8c430000; // 004008f0: LW, REG[3]<=RAM[REG[2]+0];
      10'h23d: data = 32'h8fc20008; // 004008f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h23e: data = 32'h00000000; // 004008f8: SLL, REG[0]<=REG[0]<<0;
      10'h23f: data = 32'hac430000; // 004008fc: SW, RAM[REG[2]+0]<=REG[3];
      10'h240: data = 32'h8fc20008; // 00400900: LW, REG[2]<=RAM[REG[30]+8];
      10'h241: data = 32'h00000000; // 00400904: SLL, REG[0]<=REG[0]<<0;
      10'h242: data = 32'h8c430000; // 00400908: LW, REG[3]<=RAM[REG[2]+0];
      10'h243: data = 32'h2402003e; // 0040090c: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h244: data = 32'h1462ff4f; // 00400910: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h245: data = 32'h00000000; // 00400914: SLL, REG[0]<=REG[0]<<0;
      10'h246: data = 32'h8fc20008; // 00400918: LW, REG[2]<=RAM[REG[30]+8];
      10'h247: data = 32'h00000000; // 0040091c: SLL, REG[0]<=REG[0]<<0;
      10'h248: data = 32'hac400000; // 00400920: SW, RAM[REG[2]+0]<=REG[0];
      10'h249: data = 32'h24020308; // 00400924: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h24a: data = 32'hac400000; // 00400928: SW, RAM[REG[2]+0]<=REG[0];
      10'h24b: data = 32'h2402030c; // 0040092c: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h24c: data = 32'hac400000; // 00400930: SW, RAM[REG[2]+0]<=REG[0];
      10'h24d: data = 32'h24030308; // 00400934: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h24e: data = 32'h24020001; // 00400938: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h24f: data = 32'hac620000; // 0040093c: SW, RAM[REG[3]+0]<=REG[2];
      10'h250: data = 32'h24020308; // 00400940: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h251: data = 32'hac400000; // 00400944: SW, RAM[REG[2]+0]<=REG[0];
      10'h252: data = 32'h03c0e821; // 00400948: ADDU, REG[29]<=REG[30]+REG[0];
      10'h253: data = 32'h8fbe0000; // 0040094c: LW, REG[30]<=RAM[REG[29]+0];
      10'h254: data = 32'h27bd0008; // 00400950: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h255: data = 32'h03e00008; // 00400954: JR, PC<=REG[31];
      10'h256: data = 32'h00000000; // 00400958: SLL, REG[0]<=REG[0]<<0;
      10'h257: data = 32'h27bdfff8; // 0040095c: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h258: data = 32'hafbe0000; // 00400960: SW, RAM[REG[29]+0]<=REG[30];
      10'h259: data = 32'h03a0f021; // 00400964: ADDU, REG[30]<=REG[29]+REG[0];
      10'h25a: data = 32'hafc40008; // 00400968: SW, RAM[REG[30]+8]<=REG[4];
      10'h25b: data = 32'h08100319; // 0040096c: J, PC<=0x00100319*4(=0x00400c64);
      10'h25c: data = 32'h00000000; // 00400970: SLL, REG[0]<=REG[0]<<0;
      10'h25d: data = 32'h24020300; // 00400974: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h25e: data = 32'hac400000; // 00400978: SW, RAM[REG[2]+0]<=REG[0];
      10'h25f: data = 32'h8fc20008; // 0040097c: LW, REG[2]<=RAM[REG[30]+8];
      10'h260: data = 32'h00000000; // 00400980: SLL, REG[0]<=REG[0]<<0;
      10'h261: data = 32'h8c420000; // 00400984: LW, REG[2]<=RAM[REG[2]+0];
      10'h262: data = 32'h00000000; // 00400988: SLL, REG[0]<=REG[0]<<0;
      10'h263: data = 32'h2c420041; // 0040098c: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h264: data = 32'h14400011; // 00400990: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h265: data = 32'h00000000; // 00400994: SLL, REG[0]<=REG[0]<<0;
      10'h266: data = 32'h8fc20008; // 00400998: LW, REG[2]<=RAM[REG[30]+8];
      10'h267: data = 32'h00000000; // 0040099c: SLL, REG[0]<=REG[0]<<0;
      10'h268: data = 32'h8c420000; // 004009a0: LW, REG[2]<=RAM[REG[2]+0];
      10'h269: data = 32'h00000000; // 004009a4: SLL, REG[0]<=REG[0]<<0;
      10'h26a: data = 32'h2c42005b; // 004009a8: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h26b: data = 32'h1040000a; // 004009ac: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h26c: data = 32'h00000000; // 004009b0: SLL, REG[0]<=REG[0]<<0;
      10'h26d: data = 32'h24030304; // 004009b4: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h26e: data = 32'h8fc20008; // 004009b8: LW, REG[2]<=RAM[REG[30]+8];
      10'h26f: data = 32'h00000000; // 004009bc: SLL, REG[0]<=REG[0]<<0;
      10'h270: data = 32'h8c420000; // 004009c0: LW, REG[2]<=RAM[REG[2]+0];
      10'h271: data = 32'h00000000; // 004009c4: SLL, REG[0]<=REG[0]<<0;
      10'h272: data = 32'h2442ffc0; // 004009c8: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h273: data = 32'hac620000; // 004009cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h274: data = 32'h08100312; // 004009d0: J, PC<=0x00100312*4(=0x00400c48);
      10'h275: data = 32'h00000000; // 004009d4: SLL, REG[0]<=REG[0]<<0;
      10'h276: data = 32'h8fc20008; // 004009d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h277: data = 32'h00000000; // 004009dc: SLL, REG[0]<=REG[0]<<0;
      10'h278: data = 32'h8c420000; // 004009e0: LW, REG[2]<=RAM[REG[2]+0];
      10'h279: data = 32'h00000000; // 004009e4: SLL, REG[0]<=REG[0]<<0;
      10'h27a: data = 32'h2c420061; // 004009e8: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h27b: data = 32'h14400011; // 004009ec: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h27c: data = 32'h00000000; // 004009f0: SLL, REG[0]<=REG[0]<<0;
      10'h27d: data = 32'h8fc20008; // 004009f4: LW, REG[2]<=RAM[REG[30]+8];
      10'h27e: data = 32'h00000000; // 004009f8: SLL, REG[0]<=REG[0]<<0;
      10'h27f: data = 32'h8c420000; // 004009fc: LW, REG[2]<=RAM[REG[2]+0];
      10'h280: data = 32'h00000000; // 00400a00: SLL, REG[0]<=REG[0]<<0;
      10'h281: data = 32'h2c42007b; // 00400a04: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h282: data = 32'h1040000a; // 00400a08: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h283: data = 32'h00000000; // 00400a0c: SLL, REG[0]<=REG[0]<<0;
      10'h284: data = 32'h24030304; // 00400a10: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h285: data = 32'h8fc20008; // 00400a14: LW, REG[2]<=RAM[REG[30]+8];
      10'h286: data = 32'h00000000; // 00400a18: SLL, REG[0]<=REG[0]<<0;
      10'h287: data = 32'h8c420000; // 00400a1c: LW, REG[2]<=RAM[REG[2]+0];
      10'h288: data = 32'h00000000; // 00400a20: SLL, REG[0]<=REG[0]<<0;
      10'h289: data = 32'h2442ffa0; // 00400a24: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h28a: data = 32'hac620000; // 00400a28: SW, RAM[REG[3]+0]<=REG[2];
      10'h28b: data = 32'h08100312; // 00400a2c: J, PC<=0x00100312*4(=0x00400c48);
      10'h28c: data = 32'h00000000; // 00400a30: SLL, REG[0]<=REG[0]<<0;
      10'h28d: data = 32'h8fc20008; // 00400a34: LW, REG[2]<=RAM[REG[30]+8];
      10'h28e: data = 32'h00000000; // 00400a38: SLL, REG[0]<=REG[0]<<0;
      10'h28f: data = 32'h8c420000; // 00400a3c: LW, REG[2]<=RAM[REG[2]+0];
      10'h290: data = 32'h00000000; // 00400a40: SLL, REG[0]<=REG[0]<<0;
      10'h291: data = 32'h2c420030; // 00400a44: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h292: data = 32'h14400010; // 00400a48: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h293: data = 32'h00000000; // 00400a4c: SLL, REG[0]<=REG[0]<<0;
      10'h294: data = 32'h8fc20008; // 00400a50: LW, REG[2]<=RAM[REG[30]+8];
      10'h295: data = 32'h00000000; // 00400a54: SLL, REG[0]<=REG[0]<<0;
      10'h296: data = 32'h8c420000; // 00400a58: LW, REG[2]<=RAM[REG[2]+0];
      10'h297: data = 32'h00000000; // 00400a5c: SLL, REG[0]<=REG[0]<<0;
      10'h298: data = 32'h2c42003a; // 00400a60: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h299: data = 32'h10400009; // 00400a64: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h29a: data = 32'h00000000; // 00400a68: SLL, REG[0]<=REG[0]<<0;
      10'h29b: data = 32'h24020304; // 00400a6c: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h29c: data = 32'h8fc30008; // 00400a70: LW, REG[3]<=RAM[REG[30]+8];
      10'h29d: data = 32'h00000000; // 00400a74: SLL, REG[0]<=REG[0]<<0;
      10'h29e: data = 32'h8c630000; // 00400a78: LW, REG[3]<=RAM[REG[3]+0];
      10'h29f: data = 32'h00000000; // 00400a7c: SLL, REG[0]<=REG[0]<<0;
      10'h2a0: data = 32'hac430000; // 00400a80: SW, RAM[REG[2]+0]<=REG[3];
      10'h2a1: data = 32'h08100312; // 00400a84: J, PC<=0x00100312*4(=0x00400c48);
      10'h2a2: data = 32'h00000000; // 00400a88: SLL, REG[0]<=REG[0]<<0;
      10'h2a3: data = 32'h8fc20008; // 00400a8c: LW, REG[2]<=RAM[REG[30]+8];
      10'h2a4: data = 32'h00000000; // 00400a90: SLL, REG[0]<=REG[0]<<0;
      10'h2a5: data = 32'h8c430000; // 00400a94: LW, REG[3]<=RAM[REG[2]+0];
      10'h2a6: data = 32'h24020040; // 00400a98: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h2a7: data = 32'h14620005; // 00400a9c: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h2a8: data = 32'h00000000; // 00400aa0: SLL, REG[0]<=REG[0]<<0;
      10'h2a9: data = 32'h24020304; // 00400aa4: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h2aa: data = 32'hac400000; // 00400aa8: SW, RAM[REG[2]+0]<=REG[0];
      10'h2ab: data = 32'h08100312; // 00400aac: J, PC<=0x00100312*4(=0x00400c48);
      10'h2ac: data = 32'h00000000; // 00400ab0: SLL, REG[0]<=REG[0]<<0;
      10'h2ad: data = 32'h8fc20008; // 00400ab4: LW, REG[2]<=RAM[REG[30]+8];
      10'h2ae: data = 32'h00000000; // 00400ab8: SLL, REG[0]<=REG[0]<<0;
      10'h2af: data = 32'h8c430000; // 00400abc: LW, REG[3]<=RAM[REG[2]+0];
      10'h2b0: data = 32'h2402005b; // 00400ac0: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h2b1: data = 32'h14620006; // 00400ac4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2b2: data = 32'h00000000; // 00400ac8: SLL, REG[0]<=REG[0]<<0;
      10'h2b3: data = 32'h24030304; // 00400acc: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2b4: data = 32'h2402001b; // 00400ad0: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h2b5: data = 32'hac620000; // 00400ad4: SW, RAM[REG[3]+0]<=REG[2];
      10'h2b6: data = 32'h08100312; // 00400ad8: J, PC<=0x00100312*4(=0x00400c48);
      10'h2b7: data = 32'h00000000; // 00400adc: SLL, REG[0]<=REG[0]<<0;
      10'h2b8: data = 32'h8fc20008; // 00400ae0: LW, REG[2]<=RAM[REG[30]+8];
      10'h2b9: data = 32'h00000000; // 00400ae4: SLL, REG[0]<=REG[0]<<0;
      10'h2ba: data = 32'h8c430000; // 00400ae8: LW, REG[3]<=RAM[REG[2]+0];
      10'h2bb: data = 32'h2402005d; // 00400aec: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h2bc: data = 32'h14620006; // 00400af0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2bd: data = 32'h00000000; // 00400af4: SLL, REG[0]<=REG[0]<<0;
      10'h2be: data = 32'h24030304; // 00400af8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2bf: data = 32'h2402001d; // 00400afc: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h2c0: data = 32'hac620000; // 00400b00: SW, RAM[REG[3]+0]<=REG[2];
      10'h2c1: data = 32'h08100312; // 00400b04: J, PC<=0x00100312*4(=0x00400c48);
      10'h2c2: data = 32'h00000000; // 00400b08: SLL, REG[0]<=REG[0]<<0;
      10'h2c3: data = 32'h8fc20008; // 00400b0c: LW, REG[2]<=RAM[REG[30]+8];
      10'h2c4: data = 32'h00000000; // 00400b10: SLL, REG[0]<=REG[0]<<0;
      10'h2c5: data = 32'h8c420000; // 00400b14: LW, REG[2]<=RAM[REG[2]+0];
      10'h2c6: data = 32'h00000000; // 00400b18: SLL, REG[0]<=REG[0]<<0;
      10'h2c7: data = 32'h2c420020; // 00400b1c: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h2c8: data = 32'h14400010; // 00400b20: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h2c9: data = 32'h00000000; // 00400b24: SLL, REG[0]<=REG[0]<<0;
      10'h2ca: data = 32'h8fc20008; // 00400b28: LW, REG[2]<=RAM[REG[30]+8];
      10'h2cb: data = 32'h00000000; // 00400b2c: SLL, REG[0]<=REG[0]<<0;
      10'h2cc: data = 32'h8c420000; // 00400b30: LW, REG[2]<=RAM[REG[2]+0];
      10'h2cd: data = 32'h00000000; // 00400b34: SLL, REG[0]<=REG[0]<<0;
      10'h2ce: data = 32'h2c420030; // 00400b38: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h2cf: data = 32'h10400009; // 00400b3c: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h2d0: data = 32'h00000000; // 00400b40: SLL, REG[0]<=REG[0]<<0;
      10'h2d1: data = 32'h24020304; // 00400b44: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h2d2: data = 32'h8fc30008; // 00400b48: LW, REG[3]<=RAM[REG[30]+8];
      10'h2d3: data = 32'h00000000; // 00400b4c: SLL, REG[0]<=REG[0]<<0;
      10'h2d4: data = 32'h8c630000; // 00400b50: LW, REG[3]<=RAM[REG[3]+0];
      10'h2d5: data = 32'h00000000; // 00400b54: SLL, REG[0]<=REG[0]<<0;
      10'h2d6: data = 32'hac430000; // 00400b58: SW, RAM[REG[2]+0]<=REG[3];
      10'h2d7: data = 32'h08100312; // 00400b5c: J, PC<=0x00100312*4(=0x00400c48);
      10'h2d8: data = 32'h00000000; // 00400b60: SLL, REG[0]<=REG[0]<<0;
      10'h2d9: data = 32'h8fc20008; // 00400b64: LW, REG[2]<=RAM[REG[30]+8];
      10'h2da: data = 32'h00000000; // 00400b68: SLL, REG[0]<=REG[0]<<0;
      10'h2db: data = 32'h8c430000; // 00400b6c: LW, REG[3]<=RAM[REG[2]+0];
      10'h2dc: data = 32'h2402003f; // 00400b70: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h2dd: data = 32'h14620006; // 00400b74: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2de: data = 32'h00000000; // 00400b78: SLL, REG[0]<=REG[0]<<0;
      10'h2df: data = 32'h24030304; // 00400b7c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2e0: data = 32'h2402003a; // 00400b80: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h2e1: data = 32'hac620000; // 00400b84: SW, RAM[REG[3]+0]<=REG[2];
      10'h2e2: data = 32'h08100312; // 00400b88: J, PC<=0x00100312*4(=0x00400c48);
      10'h2e3: data = 32'h00000000; // 00400b8c: SLL, REG[0]<=REG[0]<<0;
      10'h2e4: data = 32'h8fc20008; // 00400b90: LW, REG[2]<=RAM[REG[30]+8];
      10'h2e5: data = 32'h00000000; // 00400b94: SLL, REG[0]<=REG[0]<<0;
      10'h2e6: data = 32'h8c430000; // 00400b98: LW, REG[3]<=RAM[REG[2]+0];
      10'h2e7: data = 32'h2402003d; // 00400b9c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h2e8: data = 32'h14620006; // 00400ba0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2e9: data = 32'h00000000; // 00400ba4: SLL, REG[0]<=REG[0]<<0;
      10'h2ea: data = 32'h24030304; // 00400ba8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2eb: data = 32'h2402003b; // 00400bac: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h2ec: data = 32'hac620000; // 00400bb0: SW, RAM[REG[3]+0]<=REG[2];
      10'h2ed: data = 32'h08100312; // 00400bb4: J, PC<=0x00100312*4(=0x00400c48);
      10'h2ee: data = 32'h00000000; // 00400bb8: SLL, REG[0]<=REG[0]<<0;
      10'h2ef: data = 32'h8fc20008; // 00400bbc: LW, REG[2]<=RAM[REG[30]+8];
      10'h2f0: data = 32'h00000000; // 00400bc0: SLL, REG[0]<=REG[0]<<0;
      10'h2f1: data = 32'h8c430000; // 00400bc4: LW, REG[3]<=RAM[REG[2]+0];
      10'h2f2: data = 32'h2402003b; // 00400bc8: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h2f3: data = 32'h14620006; // 00400bcc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2f4: data = 32'h00000000; // 00400bd0: SLL, REG[0]<=REG[0]<<0;
      10'h2f5: data = 32'h24030304; // 00400bd4: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h2f6: data = 32'h2402003c; // 00400bd8: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h2f7: data = 32'hac620000; // 00400bdc: SW, RAM[REG[3]+0]<=REG[2];
      10'h2f8: data = 32'h08100312; // 00400be0: J, PC<=0x00100312*4(=0x00400c48);
      10'h2f9: data = 32'h00000000; // 00400be4: SLL, REG[0]<=REG[0]<<0;
      10'h2fa: data = 32'h8fc20008; // 00400be8: LW, REG[2]<=RAM[REG[30]+8];
      10'h2fb: data = 32'h00000000; // 00400bec: SLL, REG[0]<=REG[0]<<0;
      10'h2fc: data = 32'h8c430000; // 00400bf0: LW, REG[3]<=RAM[REG[2]+0];
      10'h2fd: data = 32'h2402003a; // 00400bf4: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h2fe: data = 32'h14620006; // 00400bf8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h2ff: data = 32'h00000000; // 00400bfc: SLL, REG[0]<=REG[0]<<0;
      10'h300: data = 32'h24030304; // 00400c00: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h301: data = 32'h2402003d; // 00400c04: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h302: data = 32'hac620000; // 00400c08: SW, RAM[REG[3]+0]<=REG[2];
      10'h303: data = 32'h08100312; // 00400c0c: J, PC<=0x00100312*4(=0x00400c48);
      10'h304: data = 32'h00000000; // 00400c10: SLL, REG[0]<=REG[0]<<0;
      10'h305: data = 32'h8fc20008; // 00400c14: LW, REG[2]<=RAM[REG[30]+8];
      10'h306: data = 32'h00000000; // 00400c18: SLL, REG[0]<=REG[0]<<0;
      10'h307: data = 32'h8c430000; // 00400c1c: LW, REG[3]<=RAM[REG[2]+0];
      10'h308: data = 32'h2402000a; // 00400c20: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h309: data = 32'h14620006; // 00400c24: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h30a: data = 32'h00000000; // 00400c28: SLL, REG[0]<=REG[0]<<0;
      10'h30b: data = 32'h24030304; // 00400c2c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h30c: data = 32'h2402003e; // 00400c30: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h30d: data = 32'hac620000; // 00400c34: SW, RAM[REG[3]+0]<=REG[2];
      10'h30e: data = 32'h08100312; // 00400c38: J, PC<=0x00100312*4(=0x00400c48);
      10'h30f: data = 32'h00000000; // 00400c3c: SLL, REG[0]<=REG[0]<<0;
      10'h310: data = 32'h24020304; // 00400c40: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h311: data = 32'hac400000; // 00400c44: SW, RAM[REG[2]+0]<=REG[0];
      10'h312: data = 32'h24030300; // 00400c48: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h313: data = 32'h24020001; // 00400c4c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h314: data = 32'hac620000; // 00400c50: SW, RAM[REG[3]+0]<=REG[2];
      10'h315: data = 32'h8fc20008; // 00400c54: LW, REG[2]<=RAM[REG[30]+8];
      10'h316: data = 32'h00000000; // 00400c58: SLL, REG[0]<=REG[0]<<0;
      10'h317: data = 32'h24420004; // 00400c5c: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h318: data = 32'hafc20008; // 00400c60: SW, RAM[REG[30]+8]<=REG[2];
      10'h319: data = 32'h8fc20008; // 00400c64: LW, REG[2]<=RAM[REG[30]+8];
      10'h31a: data = 32'h00000000; // 00400c68: SLL, REG[0]<=REG[0]<<0;
      10'h31b: data = 32'h8c420000; // 00400c6c: LW, REG[2]<=RAM[REG[2]+0];
      10'h31c: data = 32'h00000000; // 00400c70: SLL, REG[0]<=REG[0]<<0;
      10'h31d: data = 32'h1440ff3f; // 00400c74: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h31e: data = 32'h00000000; // 00400c78: SLL, REG[0]<=REG[0]<<0;
      10'h31f: data = 32'h03c0e821; // 00400c7c: ADDU, REG[29]<=REG[30]+REG[0];
      10'h320: data = 32'h8fbe0000; // 00400c80: LW, REG[30]<=RAM[REG[29]+0];
      10'h321: data = 32'h27bd0008; // 00400c84: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h322: data = 32'h03e00008; // 00400c88: JR, PC<=REG[31];
      10'h323: data = 32'h00000000; // 00400c8c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
