/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408740; // 00400014: SLL, REG[16]<=REG[0]<<29;
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdffa0; // 00400020: ADDIU, REG[29]<=REG[29]+65440(=0x0000ffa0);
      10'h009: data = 32'hafbf005c; // 00400024: SW, RAM[REG[29]+92]<=REG[31];
      10'h00a: data = 32'hafbe0058; // 00400028: SW, RAM[REG[29]+88]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020001; // 00400030: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h00d: data = 32'hafc20014; // 00400034: SW, RAM[REG[30]+20]<=REG[2];
      10'h00e: data = 32'h27c20018; // 00400038: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h00f: data = 32'h00402021; // 0040003c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h010: data = 32'h0c10005c; // 00400040: JAL, PC<=0x0010005c*4(=0x00400170); REG[31]<=PC+4
      10'h011: data = 32'h00000000; // 00400044: SLL, REG[0]<=REG[0]<<0;
      10'h012: data = 32'h27c20018; // 00400048: ADDIU, REG[2]<=REG[30]+24(=0x00000018);
      10'h013: data = 32'h00402021; // 0040004c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h014: data = 32'h0c10013e; // 00400050: JAL, PC<=0x0010013e*4(=0x004004f8); REG[31]<=PC+4
      10'h015: data = 32'h00000000; // 00400054: SLL, REG[0]<=REG[0]<<0;
      10'h016: data = 32'hafc20010; // 00400058: SW, RAM[REG[30]+16]<=REG[2];
      10'h017: data = 32'h8fc30010; // 0040005c: LW, REG[3]<=RAM[REG[30]+16];
      10'h018: data = 32'h24020002; // 00400060: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h019: data = 32'h14620005; // 00400064: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h01a: data = 32'h00000000; // 00400068: SLL, REG[0]<=REG[0]<<0;
      10'h01b: data = 32'h0c100039; // 0040006c: JAL, PC<=0x00100039*4(=0x004000e4); REG[31]<=PC+4
      10'h01c: data = 32'h00000000; // 00400070: SLL, REG[0]<=REG[0]<<0;
      10'h01d: data = 32'h08100017; // 00400074: J, PC<=0x00100017*4(=0x0040005c);
      10'h01e: data = 32'h00000000; // 00400078: SLL, REG[0]<=REG[0]<<0;
      10'h01f: data = 32'h0c100023; // 0040007c: JAL, PC<=0x00100023*4(=0x0040008c); REG[31]<=PC+4
      10'h020: data = 32'h00000000; // 00400080: SLL, REG[0]<=REG[0]<<0;
      10'h021: data = 32'h08100017; // 00400084: J, PC<=0x00100017*4(=0x0040005c);
      10'h022: data = 32'h00000000; // 00400088: SLL, REG[0]<=REG[0]<<0;
      10'h023: data = 32'h27bdffe8; // 0040008c: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h024: data = 32'hafbf0014; // 00400090: SW, RAM[REG[29]+20]<=REG[31];
      10'h025: data = 32'hafbe0010; // 00400094: SW, RAM[REG[29]+16]<=REG[30];
      10'h026: data = 32'h03a0f021; // 00400098: ADDU, REG[30]<=REG[29]+REG[0];
      10'h027: data = 32'h24040008; // 0040009c: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h028: data = 32'h0c10004f; // 004000a0: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h029: data = 32'h00000000; // 004000a4: SLL, REG[0]<=REG[0]<<0;
      10'h02a: data = 32'h24040004; // 004000a8: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h02b: data = 32'h0c10004f; // 004000ac: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h02c: data = 32'h00000000; // 004000b0: SLL, REG[0]<=REG[0]<<0;
      10'h02d: data = 32'h24040002; // 004000b4: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h02e: data = 32'h0c10004f; // 004000b8: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h02f: data = 32'h00000000; // 004000bc: SLL, REG[0]<=REG[0]<<0;
      10'h030: data = 32'h24040001; // 004000c0: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h031: data = 32'h0c10004f; // 004000c4: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h032: data = 32'h00000000; // 004000c8: SLL, REG[0]<=REG[0]<<0;
      10'h033: data = 32'h03c0e821; // 004000cc: ADDU, REG[29]<=REG[30]+REG[0];
      10'h034: data = 32'h8fbf0014; // 004000d0: LW, REG[31]<=RAM[REG[29]+20];
      10'h035: data = 32'h8fbe0010; // 004000d4: LW, REG[30]<=RAM[REG[29]+16];
      10'h036: data = 32'h27bd0018; // 004000d8: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h037: data = 32'h03e00008; // 004000dc: JR, PC<=REG[31];
      10'h038: data = 32'h00000000; // 004000e0: SLL, REG[0]<=REG[0]<<0;
      10'h039: data = 32'h27bdffe8; // 004000e4: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h03a: data = 32'hafbf0014; // 004000e8: SW, RAM[REG[29]+20]<=REG[31];
      10'h03b: data = 32'hafbe0010; // 004000ec: SW, RAM[REG[29]+16]<=REG[30];
      10'h03c: data = 32'h03a0f021; // 004000f0: ADDU, REG[30]<=REG[29]+REG[0];
      10'h03d: data = 32'h24040001; // 004000f4: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h03e: data = 32'h0c10004f; // 004000f8: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h03f: data = 32'h00000000; // 004000fc: SLL, REG[0]<=REG[0]<<0;
      10'h040: data = 32'h24040002; // 00400100: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h041: data = 32'h0c10004f; // 00400104: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h042: data = 32'h00000000; // 00400108: SLL, REG[0]<=REG[0]<<0;
      10'h043: data = 32'h24040004; // 0040010c: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h044: data = 32'h0c10004f; // 00400110: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h045: data = 32'h00000000; // 00400114: SLL, REG[0]<=REG[0]<<0;
      10'h046: data = 32'h24040008; // 00400118: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h047: data = 32'h0c10004f; // 0040011c: JAL, PC<=0x0010004f*4(=0x0040013c); REG[31]<=PC+4
      10'h048: data = 32'h00000000; // 00400120: SLL, REG[0]<=REG[0]<<0;
      10'h049: data = 32'h03c0e821; // 00400124: ADDU, REG[29]<=REG[30]+REG[0];
      10'h04a: data = 32'h8fbf0014; // 00400128: LW, REG[31]<=RAM[REG[29]+20];
      10'h04b: data = 32'h8fbe0010; // 0040012c: LW, REG[30]<=RAM[REG[29]+16];
      10'h04c: data = 32'h27bd0018; // 00400130: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h04d: data = 32'h03e00008; // 00400134: JR, PC<=REG[31];
      10'h04e: data = 32'h00000000; // 00400138: SLL, REG[0]<=REG[0]<<0;
      10'h04f: data = 32'h27bdfff0; // 0040013c: ADDIU, REG[29]<=REG[29]+65520(=0x0000fff0);
      10'h050: data = 32'hafbe0008; // 00400140: SW, RAM[REG[29]+8]<=REG[30];
      10'h051: data = 32'h03a0f021; // 00400144: ADDU, REG[30]<=REG[29]+REG[0];
      10'h052: data = 32'hafc40010; // 00400148: SW, RAM[REG[30]+16]<=REG[4];
      10'h053: data = 32'h24030320; // 0040014c: ADDIU, REG[3]<=REG[0]+800(=0x00000320);
      10'h054: data = 32'h8fc20010; // 00400150: LW, REG[2]<=RAM[REG[30]+16];
      10'h055: data = 32'h00000000; // 00400154: SLL, REG[0]<=REG[0]<<0;
      10'h056: data = 32'hac620000; // 00400158: SW, RAM[REG[3]+0]<=REG[2];
      10'h057: data = 32'h03c0e821; // 0040015c: ADDU, REG[29]<=REG[30]+REG[0];
      10'h058: data = 32'h8fbe0008; // 00400160: LW, REG[30]<=RAM[REG[29]+8];
      10'h059: data = 32'h27bd0010; // 00400164: ADDIU, REG[29]<=REG[29]+16(=0x00000010);
      10'h05a: data = 32'h03e00008; // 00400168: JR, PC<=REG[31];
      10'h05b: data = 32'h00000000; // 0040016c: SLL, REG[0]<=REG[0]<<0;
      10'h05c: data = 32'h27bdfff8; // 00400170: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h05d: data = 32'hafbe0000; // 00400174: SW, RAM[REG[29]+0]<=REG[30];
      10'h05e: data = 32'h03a0f021; // 00400178: ADDU, REG[30]<=REG[29]+REG[0];
      10'h05f: data = 32'hafc40008; // 0040017c: SW, RAM[REG[30]+8]<=REG[4];
      10'h060: data = 32'h24020308; // 00400180: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h061: data = 32'hac400000; // 00400184: SW, RAM[REG[2]+0]<=REG[0];
      10'h062: data = 32'h2403030c; // 00400188: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h063: data = 32'h24020001; // 0040018c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h064: data = 32'hac620000; // 00400190: SW, RAM[REG[3]+0]<=REG[2];
      10'h065: data = 32'h24030308; // 00400194: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h066: data = 32'h24020001; // 00400198: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h067: data = 32'hac620000; // 0040019c: SW, RAM[REG[3]+0]<=REG[2];
      10'h068: data = 32'h24020308; // 004001a0: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h069: data = 32'hac400000; // 004001a4: SW, RAM[REG[2]+0]<=REG[0];
      10'h06a: data = 32'h24030308; // 004001a8: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h06b: data = 32'h24020001; // 004001ac: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h06c: data = 32'hac620000; // 004001b0: SW, RAM[REG[3]+0]<=REG[2];
      10'h06d: data = 32'h08100074; // 004001b4: J, PC<=0x00100074*4(=0x004001d0);
      10'h06e: data = 32'h00000000; // 004001b8: SLL, REG[0]<=REG[0]<<0;
      10'h06f: data = 32'h24020308; // 004001bc: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h070: data = 32'hac400000; // 004001c0: SW, RAM[REG[2]+0]<=REG[0];
      10'h071: data = 32'h24030308; // 004001c4: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h072: data = 32'h24020001; // 004001c8: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h073: data = 32'hac620000; // 004001cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h074: data = 32'h24020310; // 004001d0: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h075: data = 32'h8c430000; // 004001d4: LW, REG[3]<=RAM[REG[2]+0];
      10'h076: data = 32'h2402ffff; // 004001d8: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h077: data = 32'h1062fff7; // 004001dc: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h078: data = 32'h00000000; // 004001e0: SLL, REG[0]<=REG[0]<<0;
      10'h079: data = 32'h08100122; // 004001e4: J, PC<=0x00100122*4(=0x00400488);
      10'h07a: data = 32'h00000000; // 004001e8: SLL, REG[0]<=REG[0]<<0;
      10'h07b: data = 32'h8fc20008; // 004001ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h07c: data = 32'h00000000; // 004001f0: SLL, REG[0]<=REG[0]<<0;
      10'h07d: data = 32'h8c420000; // 004001f4: LW, REG[2]<=RAM[REG[2]+0];
      10'h07e: data = 32'h00000000; // 004001f8: SLL, REG[0]<=REG[0]<<0;
      10'h07f: data = 32'h10400012; // 004001fc: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h080: data = 32'h00000000; // 00400200: SLL, REG[0]<=REG[0]<<0;
      10'h081: data = 32'h8fc20008; // 00400204: LW, REG[2]<=RAM[REG[30]+8];
      10'h082: data = 32'h00000000; // 00400208: SLL, REG[0]<=REG[0]<<0;
      10'h083: data = 32'h8c420000; // 0040020c: LW, REG[2]<=RAM[REG[2]+0];
      10'h084: data = 32'h00000000; // 00400210: SLL, REG[0]<=REG[0]<<0;
      10'h085: data = 32'h2c42001b; // 00400214: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h086: data = 32'h1040000b; // 00400218: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h087: data = 32'h00000000; // 0040021c: SLL, REG[0]<=REG[0]<<0;
      10'h088: data = 32'h8fc20008; // 00400220: LW, REG[2]<=RAM[REG[30]+8];
      10'h089: data = 32'h00000000; // 00400224: SLL, REG[0]<=REG[0]<<0;
      10'h08a: data = 32'h8c420000; // 00400228: LW, REG[2]<=RAM[REG[2]+0];
      10'h08b: data = 32'h00000000; // 0040022c: SLL, REG[0]<=REG[0]<<0;
      10'h08c: data = 32'h24430040; // 00400230: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h08d: data = 32'h8fc20008; // 00400234: LW, REG[2]<=RAM[REG[30]+8];
      10'h08e: data = 32'h00000000; // 00400238: SLL, REG[0]<=REG[0]<<0;
      10'h08f: data = 32'hac430000; // 0040023c: SW, RAM[REG[2]+0]<=REG[3];
      10'h090: data = 32'h08100119; // 00400240: J, PC<=0x00100119*4(=0x00400464);
      10'h091: data = 32'h00000000; // 00400244: SLL, REG[0]<=REG[0]<<0;
      10'h092: data = 32'h8fc20008; // 00400248: LW, REG[2]<=RAM[REG[30]+8];
      10'h093: data = 32'h00000000; // 0040024c: SLL, REG[0]<=REG[0]<<0;
      10'h094: data = 32'h8c420000; // 00400250: LW, REG[2]<=RAM[REG[2]+0];
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h2c420030; // 00400258: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h097: data = 32'h14400010; // 0040025c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h098: data = 32'h00000000; // 00400260: SLL, REG[0]<=REG[0]<<0;
      10'h099: data = 32'h8fc20008; // 00400264: LW, REG[2]<=RAM[REG[30]+8];
      10'h09a: data = 32'h00000000; // 00400268: SLL, REG[0]<=REG[0]<<0;
      10'h09b: data = 32'h8c420000; // 0040026c: LW, REG[2]<=RAM[REG[2]+0];
      10'h09c: data = 32'h00000000; // 00400270: SLL, REG[0]<=REG[0]<<0;
      10'h09d: data = 32'h2c42003a; // 00400274: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h09e: data = 32'h10400009; // 00400278: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h09f: data = 32'h00000000; // 0040027c: SLL, REG[0]<=REG[0]<<0;
      10'h0a0: data = 32'h8fc20008; // 00400280: LW, REG[2]<=RAM[REG[30]+8];
      10'h0a1: data = 32'h00000000; // 00400284: SLL, REG[0]<=REG[0]<<0;
      10'h0a2: data = 32'h8c430000; // 00400288: LW, REG[3]<=RAM[REG[2]+0];
      10'h0a3: data = 32'h8fc20008; // 0040028c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0a4: data = 32'h00000000; // 00400290: SLL, REG[0]<=REG[0]<<0;
      10'h0a5: data = 32'hac430000; // 00400294: SW, RAM[REG[2]+0]<=REG[3];
      10'h0a6: data = 32'h08100119; // 00400298: J, PC<=0x00100119*4(=0x00400464);
      10'h0a7: data = 32'h00000000; // 0040029c: SLL, REG[0]<=REG[0]<<0;
      10'h0a8: data = 32'h8fc20008; // 004002a0: LW, REG[2]<=RAM[REG[30]+8];
      10'h0a9: data = 32'h00000000; // 004002a4: SLL, REG[0]<=REG[0]<<0;
      10'h0aa: data = 32'h8c420000; // 004002a8: LW, REG[2]<=RAM[REG[2]+0];
      10'h0ab: data = 32'h00000000; // 004002ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ac: data = 32'h14400006; // 004002b0: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h0ad: data = 32'h00000000; // 004002b4: SLL, REG[0]<=REG[0]<<0;
      10'h0ae: data = 32'h8fc30008; // 004002b8: LW, REG[3]<=RAM[REG[30]+8];
      10'h0af: data = 32'h24020040; // 004002bc: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h0b0: data = 32'hac620000; // 004002c0: SW, RAM[REG[3]+0]<=REG[2];
      10'h0b1: data = 32'h08100119; // 004002c4: J, PC<=0x00100119*4(=0x00400464);
      10'h0b2: data = 32'h00000000; // 004002c8: SLL, REG[0]<=REG[0]<<0;
      10'h0b3: data = 32'h8fc20008; // 004002cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b4: data = 32'h00000000; // 004002d0: SLL, REG[0]<=REG[0]<<0;
      10'h0b5: data = 32'h8c430000; // 004002d4: LW, REG[3]<=RAM[REG[2]+0];
      10'h0b6: data = 32'h2402001b; // 004002d8: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h0b7: data = 32'h14620006; // 004002dc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0b8: data = 32'h00000000; // 004002e0: SLL, REG[0]<=REG[0]<<0;
      10'h0b9: data = 32'h8fc30008; // 004002e4: LW, REG[3]<=RAM[REG[30]+8];
      10'h0ba: data = 32'h2402005b; // 004002e8: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h0bb: data = 32'hac620000; // 004002ec: SW, RAM[REG[3]+0]<=REG[2];
      10'h0bc: data = 32'h08100119; // 004002f0: J, PC<=0x00100119*4(=0x00400464);
      10'h0bd: data = 32'h00000000; // 004002f4: SLL, REG[0]<=REG[0]<<0;
      10'h0be: data = 32'h8fc20008; // 004002f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0bf: data = 32'h00000000; // 004002fc: SLL, REG[0]<=REG[0]<<0;
      10'h0c0: data = 32'h8c430000; // 00400300: LW, REG[3]<=RAM[REG[2]+0];
      10'h0c1: data = 32'h2402001d; // 00400304: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h0c2: data = 32'h14620006; // 00400308: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0c3: data = 32'h00000000; // 0040030c: SLL, REG[0]<=REG[0]<<0;
      10'h0c4: data = 32'h8fc30008; // 00400310: LW, REG[3]<=RAM[REG[30]+8];
      10'h0c5: data = 32'h2402005d; // 00400314: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h0c6: data = 32'hac620000; // 00400318: SW, RAM[REG[3]+0]<=REG[2];
      10'h0c7: data = 32'h08100119; // 0040031c: J, PC<=0x00100119*4(=0x00400464);
      10'h0c8: data = 32'h00000000; // 00400320: SLL, REG[0]<=REG[0]<<0;
      10'h0c9: data = 32'h8fc20008; // 00400324: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ca: data = 32'h00000000; // 00400328: SLL, REG[0]<=REG[0]<<0;
      10'h0cb: data = 32'h8c420000; // 0040032c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cc: data = 32'h00000000; // 00400330: SLL, REG[0]<=REG[0]<<0;
      10'h0cd: data = 32'h2c420020; // 00400334: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h0ce: data = 32'h14400010; // 00400338: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h0cf: data = 32'h00000000; // 0040033c: SLL, REG[0]<=REG[0]<<0;
      10'h0d0: data = 32'h8fc20008; // 00400340: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d1: data = 32'h00000000; // 00400344: SLL, REG[0]<=REG[0]<<0;
      10'h0d2: data = 32'h8c420000; // 00400348: LW, REG[2]<=RAM[REG[2]+0];
      10'h0d3: data = 32'h00000000; // 0040034c: SLL, REG[0]<=REG[0]<<0;
      10'h0d4: data = 32'h2c420030; // 00400350: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0d5: data = 32'h10400009; // 00400354: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0d6: data = 32'h00000000; // 00400358: SLL, REG[0]<=REG[0]<<0;
      10'h0d7: data = 32'h8fc20008; // 0040035c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d8: data = 32'h00000000; // 00400360: SLL, REG[0]<=REG[0]<<0;
      10'h0d9: data = 32'h8c430000; // 00400364: LW, REG[3]<=RAM[REG[2]+0];
      10'h0da: data = 32'h8fc20008; // 00400368: LW, REG[2]<=RAM[REG[30]+8];
      10'h0db: data = 32'h00000000; // 0040036c: SLL, REG[0]<=REG[0]<<0;
      10'h0dc: data = 32'hac430000; // 00400370: SW, RAM[REG[2]+0]<=REG[3];
      10'h0dd: data = 32'h08100119; // 00400374: J, PC<=0x00100119*4(=0x00400464);
      10'h0de: data = 32'h00000000; // 00400378: SLL, REG[0]<=REG[0]<<0;
      10'h0df: data = 32'h8fc20008; // 0040037c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e0: data = 32'h00000000; // 00400380: SLL, REG[0]<=REG[0]<<0;
      10'h0e1: data = 32'h8c430000; // 00400384: LW, REG[3]<=RAM[REG[2]+0];
      10'h0e2: data = 32'h2402003a; // 00400388: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h0e3: data = 32'h14620006; // 0040038c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0e4: data = 32'h00000000; // 00400390: SLL, REG[0]<=REG[0]<<0;
      10'h0e5: data = 32'h8fc30008; // 00400394: LW, REG[3]<=RAM[REG[30]+8];
      10'h0e6: data = 32'h2402003f; // 00400398: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h0e7: data = 32'hac620000; // 0040039c: SW, RAM[REG[3]+0]<=REG[2];
      10'h0e8: data = 32'h08100119; // 004003a0: J, PC<=0x00100119*4(=0x00400464);
      10'h0e9: data = 32'h00000000; // 004003a4: SLL, REG[0]<=REG[0]<<0;
      10'h0ea: data = 32'h8fc20008; // 004003a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0eb: data = 32'h00000000; // 004003ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ec: data = 32'h8c430000; // 004003b0: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ed: data = 32'h2402003b; // 004003b4: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0ee: data = 32'h14620006; // 004003b8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0ef: data = 32'h00000000; // 004003bc: SLL, REG[0]<=REG[0]<<0;
      10'h0f0: data = 32'h8fc30008; // 004003c0: LW, REG[3]<=RAM[REG[30]+8];
      10'h0f1: data = 32'h2402003d; // 004003c4: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h0f2: data = 32'hac620000; // 004003c8: SW, RAM[REG[3]+0]<=REG[2];
      10'h0f3: data = 32'h08100119; // 004003cc: J, PC<=0x00100119*4(=0x00400464);
      10'h0f4: data = 32'h00000000; // 004003d0: SLL, REG[0]<=REG[0]<<0;
      10'h0f5: data = 32'h8fc20008; // 004003d4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f6: data = 32'h00000000; // 004003d8: SLL, REG[0]<=REG[0]<<0;
      10'h0f7: data = 32'h8c430000; // 004003dc: LW, REG[3]<=RAM[REG[2]+0];
      10'h0f8: data = 32'h2402003c; // 004003e0: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h0f9: data = 32'h14620006; // 004003e4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0fa: data = 32'h00000000; // 004003e8: SLL, REG[0]<=REG[0]<<0;
      10'h0fb: data = 32'h8fc30008; // 004003ec: LW, REG[3]<=RAM[REG[30]+8];
      10'h0fc: data = 32'h2402003b; // 004003f0: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h0fd: data = 32'hac620000; // 004003f4: SW, RAM[REG[3]+0]<=REG[2];
      10'h0fe: data = 32'h08100119; // 004003f8: J, PC<=0x00100119*4(=0x00400464);
      10'h0ff: data = 32'h00000000; // 004003fc: SLL, REG[0]<=REG[0]<<0;
      10'h100: data = 32'h8fc20008; // 00400400: LW, REG[2]<=RAM[REG[30]+8];
      10'h101: data = 32'h00000000; // 00400404: SLL, REG[0]<=REG[0]<<0;
      10'h102: data = 32'h8c430000; // 00400408: LW, REG[3]<=RAM[REG[2]+0];
      10'h103: data = 32'h2402003d; // 0040040c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h104: data = 32'h14620006; // 00400410: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h105: data = 32'h00000000; // 00400414: SLL, REG[0]<=REG[0]<<0;
      10'h106: data = 32'h8fc30008; // 00400418: LW, REG[3]<=RAM[REG[30]+8];
      10'h107: data = 32'h2402003a; // 0040041c: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h108: data = 32'hac620000; // 00400420: SW, RAM[REG[3]+0]<=REG[2];
      10'h109: data = 32'h08100119; // 00400424: J, PC<=0x00100119*4(=0x00400464);
      10'h10a: data = 32'h00000000; // 00400428: SLL, REG[0]<=REG[0]<<0;
      10'h10b: data = 32'h8fc20008; // 0040042c: LW, REG[2]<=RAM[REG[30]+8];
      10'h10c: data = 32'h00000000; // 00400430: SLL, REG[0]<=REG[0]<<0;
      10'h10d: data = 32'h8c430000; // 00400434: LW, REG[3]<=RAM[REG[2]+0];
      10'h10e: data = 32'h2402003e; // 00400438: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h10f: data = 32'h14620006; // 0040043c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h110: data = 32'h00000000; // 00400440: SLL, REG[0]<=REG[0]<<0;
      10'h111: data = 32'h8fc30008; // 00400444: LW, REG[3]<=RAM[REG[30]+8];
      10'h112: data = 32'h2402000a; // 00400448: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h113: data = 32'hac620000; // 0040044c: SW, RAM[REG[3]+0]<=REG[2];
      10'h114: data = 32'h08100119; // 00400450: J, PC<=0x00100119*4(=0x00400464);
      10'h115: data = 32'h00000000; // 00400454: SLL, REG[0]<=REG[0]<<0;
      10'h116: data = 32'h8fc30008; // 00400458: LW, REG[3]<=RAM[REG[30]+8];
      10'h117: data = 32'h24020040; // 0040045c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h118: data = 32'hac620000; // 00400460: SW, RAM[REG[3]+0]<=REG[2];
      10'h119: data = 32'h24020308; // 00400464: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h11a: data = 32'hac400000; // 00400468: SW, RAM[REG[2]+0]<=REG[0];
      10'h11b: data = 32'h24030308; // 0040046c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h11c: data = 32'h24020001; // 00400470: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h11d: data = 32'hac620000; // 00400474: SW, RAM[REG[3]+0]<=REG[2];
      10'h11e: data = 32'h8fc20008; // 00400478: LW, REG[2]<=RAM[REG[30]+8];
      10'h11f: data = 32'h00000000; // 0040047c: SLL, REG[0]<=REG[0]<<0;
      10'h120: data = 32'h24420004; // 00400480: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h121: data = 32'hafc20008; // 00400484: SW, RAM[REG[30]+8]<=REG[2];
      10'h122: data = 32'h24020310; // 00400488: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h123: data = 32'h8c430000; // 0040048c: LW, REG[3]<=RAM[REG[2]+0];
      10'h124: data = 32'h8fc20008; // 00400490: LW, REG[2]<=RAM[REG[30]+8];
      10'h125: data = 32'h00000000; // 00400494: SLL, REG[0]<=REG[0]<<0;
      10'h126: data = 32'hac430000; // 00400498: SW, RAM[REG[2]+0]<=REG[3];
      10'h127: data = 32'h8fc20008; // 0040049c: LW, REG[2]<=RAM[REG[30]+8];
      10'h128: data = 32'h00000000; // 004004a0: SLL, REG[0]<=REG[0]<<0;
      10'h129: data = 32'h8c430000; // 004004a4: LW, REG[3]<=RAM[REG[2]+0];
      10'h12a: data = 32'h2402003e; // 004004a8: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h12b: data = 32'h1462ff4f; // 004004ac: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h12c: data = 32'h00000000; // 004004b0: SLL, REG[0]<=REG[0]<<0;
      10'h12d: data = 32'h8fc20008; // 004004b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h12e: data = 32'h00000000; // 004004b8: SLL, REG[0]<=REG[0]<<0;
      10'h12f: data = 32'hac400000; // 004004bc: SW, RAM[REG[2]+0]<=REG[0];
      10'h130: data = 32'h24020308; // 004004c0: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h131: data = 32'hac400000; // 004004c4: SW, RAM[REG[2]+0]<=REG[0];
      10'h132: data = 32'h2402030c; // 004004c8: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h133: data = 32'hac400000; // 004004cc: SW, RAM[REG[2]+0]<=REG[0];
      10'h134: data = 32'h24030308; // 004004d0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h135: data = 32'h24020001; // 004004d4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h136: data = 32'hac620000; // 004004d8: SW, RAM[REG[3]+0]<=REG[2];
      10'h137: data = 32'h24020308; // 004004dc: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h138: data = 32'hac400000; // 004004e0: SW, RAM[REG[2]+0]<=REG[0];
      10'h139: data = 32'h03c0e821; // 004004e4: ADDU, REG[29]<=REG[30]+REG[0];
      10'h13a: data = 32'h8fbe0000; // 004004e8: LW, REG[30]<=RAM[REG[29]+0];
      10'h13b: data = 32'h27bd0008; // 004004ec: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h13c: data = 32'h03e00008; // 004004f0: JR, PC<=REG[31];
      10'h13d: data = 32'h00000000; // 004004f4: SLL, REG[0]<=REG[0]<<0;
      10'h13e: data = 32'h27bdffe8; // 004004f8: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h13f: data = 32'hafbe0010; // 004004fc: SW, RAM[REG[29]+16]<=REG[30];
      10'h140: data = 32'h03a0f021; // 00400500: ADDU, REG[30]<=REG[29]+REG[0];
      10'h141: data = 32'hafc40018; // 00400504: SW, RAM[REG[30]+24]<=REG[4];
      10'h142: data = 32'h8fc20018; // 00400508: LW, REG[2]<=RAM[REG[30]+24];
      10'h143: data = 32'h00000000; // 0040050c: SLL, REG[0]<=REG[0]<<0;
      10'h144: data = 32'hafc20008; // 00400510: SW, RAM[REG[30]+8]<=REG[2];
      10'h145: data = 32'hafc00004; // 00400514: SW, RAM[REG[30]+4]<=REG[0];
      10'h146: data = 32'h08100150; // 00400518: J, PC<=0x00100150*4(=0x00400540);
      10'h147: data = 32'h00000000; // 0040051c: SLL, REG[0]<=REG[0]<<0;
      10'h148: data = 32'h8fc20008; // 00400520: LW, REG[2]<=RAM[REG[30]+8];
      10'h149: data = 32'h00000000; // 00400524: SLL, REG[0]<=REG[0]<<0;
      10'h14a: data = 32'h24420004; // 00400528: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h14b: data = 32'hafc20008; // 0040052c: SW, RAM[REG[30]+8]<=REG[2];
      10'h14c: data = 32'h8fc20004; // 00400530: LW, REG[2]<=RAM[REG[30]+4];
      10'h14d: data = 32'h00000000; // 00400534: SLL, REG[0]<=REG[0]<<0;
      10'h14e: data = 32'h24420001; // 00400538: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h14f: data = 32'hafc20004; // 0040053c: SW, RAM[REG[30]+4]<=REG[2];
      10'h150: data = 32'h8fc20008; // 00400540: LW, REG[2]<=RAM[REG[30]+8];
      10'h151: data = 32'h00000000; // 00400544: SLL, REG[0]<=REG[0]<<0;
      10'h152: data = 32'h8c420000; // 00400548: LW, REG[2]<=RAM[REG[2]+0];
      10'h153: data = 32'h00000000; // 0040054c: SLL, REG[0]<=REG[0]<<0;
      10'h154: data = 32'h1440fff3; // 00400550: BNE, PC<=(REG[2] != REG[0])?PC+4+65523*4:PC+4;
      10'h155: data = 32'h00000000; // 00400554: SLL, REG[0]<=REG[0]<<0;
      10'h156: data = 32'hafc00000; // 00400558: SW, RAM[REG[30]+0]<=REG[0];
      10'h157: data = 32'h8fc20018; // 0040055c: LW, REG[2]<=RAM[REG[30]+24];
      10'h158: data = 32'h00000000; // 00400560: SLL, REG[0]<=REG[0]<<0;
      10'h159: data = 32'hafc20008; // 00400564: SW, RAM[REG[30]+8]<=REG[2];
      10'h15a: data = 32'h8fc30004; // 00400568: LW, REG[3]<=RAM[REG[30]+4];
      10'h15b: data = 32'h24020001; // 0040056c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h15c: data = 32'h14620009; // 00400570: BNE, PC<=(REG[3] != REG[2])?PC+4+9*4:PC+4;
      10'h15d: data = 32'h00000000; // 00400574: SLL, REG[0]<=REG[0]<<0;
      10'h15e: data = 32'h8fc20008; // 00400578: LW, REG[2]<=RAM[REG[30]+8];
      10'h15f: data = 32'h00000000; // 0040057c: SLL, REG[0]<=REG[0]<<0;
      10'h160: data = 32'h8c420000; // 00400580: LW, REG[2]<=RAM[REG[2]+0];
      10'h161: data = 32'h00000000; // 00400584: SLL, REG[0]<=REG[0]<<0;
      10'h162: data = 32'h2442ffd0; // 00400588: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h163: data = 32'hafc20000; // 0040058c: SW, RAM[REG[30]+0]<=REG[2];
      10'h164: data = 32'h081001cb; // 00400590: J, PC<=0x001001cb*4(=0x0040072c);
      10'h165: data = 32'h00000000; // 00400594: SLL, REG[0]<=REG[0]<<0;
      10'h166: data = 32'h8fc30004; // 00400598: LW, REG[3]<=RAM[REG[30]+4];
      10'h167: data = 32'h24020002; // 0040059c: ADDIU, REG[2]<=REG[0]+2(=0x00000002);
      10'h168: data = 32'h14620024; // 004005a0: BNE, PC<=(REG[3] != REG[2])?PC+4+36*4:PC+4;
      10'h169: data = 32'h00000000; // 004005a4: SLL, REG[0]<=REG[0]<<0;
      10'h16a: data = 32'hafc00004; // 004005a8: SW, RAM[REG[30]+4]<=REG[0];
      10'h16b: data = 32'h08100175; // 004005ac: J, PC<=0x00100175*4(=0x004005d4);
      10'h16c: data = 32'h00000000; // 004005b0: SLL, REG[0]<=REG[0]<<0;
      10'h16d: data = 32'h8fc20000; // 004005b4: LW, REG[2]<=RAM[REG[30]+0];
      10'h16e: data = 32'h00000000; // 004005b8: SLL, REG[0]<=REG[0]<<0;
      10'h16f: data = 32'h2442000a; // 004005bc: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h170: data = 32'hafc20000; // 004005c0: SW, RAM[REG[30]+0]<=REG[2];
      10'h171: data = 32'h8fc20004; // 004005c4: LW, REG[2]<=RAM[REG[30]+4];
      10'h172: data = 32'h00000000; // 004005c8: SLL, REG[0]<=REG[0]<<0;
      10'h173: data = 32'h24420001; // 004005cc: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h174: data = 32'hafc20004; // 004005d0: SW, RAM[REG[30]+4]<=REG[2];
      10'h175: data = 32'h8fc20008; // 004005d4: LW, REG[2]<=RAM[REG[30]+8];
      10'h176: data = 32'h00000000; // 004005d8: SLL, REG[0]<=REG[0]<<0;
      10'h177: data = 32'h8c420000; // 004005dc: LW, REG[2]<=RAM[REG[2]+0];
      10'h178: data = 32'h00000000; // 004005e0: SLL, REG[0]<=REG[0]<<0;
      10'h179: data = 32'h2443ffd0; // 004005e4: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h17a: data = 32'h8fc20004; // 004005e8: LW, REG[2]<=RAM[REG[30]+4];
      10'h17b: data = 32'h00000000; // 004005ec: SLL, REG[0]<=REG[0]<<0;
      10'h17c: data = 32'h0043102b; // 004005f0: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h17d: data = 32'h1440ffef; // 004005f4: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h17e: data = 32'h00000000; // 004005f8: SLL, REG[0]<=REG[0]<<0;
      10'h17f: data = 32'h8fc20008; // 004005fc: LW, REG[2]<=RAM[REG[30]+8];
      10'h180: data = 32'h00000000; // 00400600: SLL, REG[0]<=REG[0]<<0;
      10'h181: data = 32'h24420004; // 00400604: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h182: data = 32'hafc20008; // 00400608: SW, RAM[REG[30]+8]<=REG[2];
      10'h183: data = 32'h8fc20008; // 0040060c: LW, REG[2]<=RAM[REG[30]+8];
      10'h184: data = 32'h00000000; // 00400610: SLL, REG[0]<=REG[0]<<0;
      10'h185: data = 32'h8c430000; // 00400614: LW, REG[3]<=RAM[REG[2]+0];
      10'h186: data = 32'h8fc20000; // 00400618: LW, REG[2]<=RAM[REG[30]+0];
      10'h187: data = 32'h00000000; // 0040061c: SLL, REG[0]<=REG[0]<<0;
      10'h188: data = 32'h00621021; // 00400620: ADDU, REG[2]<=REG[3]+REG[2];
      10'h189: data = 32'h2442ffd0; // 00400624: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h18a: data = 32'hafc20000; // 00400628: SW, RAM[REG[30]+0]<=REG[2];
      10'h18b: data = 32'h081001cb; // 0040062c: J, PC<=0x001001cb*4(=0x0040072c);
      10'h18c: data = 32'h00000000; // 00400630: SLL, REG[0]<=REG[0]<<0;
      10'h18d: data = 32'h8fc30004; // 00400634: LW, REG[3]<=RAM[REG[30]+4];
      10'h18e: data = 32'h24020003; // 00400638: ADDIU, REG[2]<=REG[0]+3(=0x00000003);
      10'h18f: data = 32'h1462003b; // 0040063c: BNE, PC<=(REG[3] != REG[2])?PC+4+59*4:PC+4;
      10'h190: data = 32'h00000000; // 00400640: SLL, REG[0]<=REG[0]<<0;
      10'h191: data = 32'hafc00004; // 00400644: SW, RAM[REG[30]+4]<=REG[0];
      10'h192: data = 32'h0810019c; // 00400648: J, PC<=0x0010019c*4(=0x00400670);
      10'h193: data = 32'h00000000; // 0040064c: SLL, REG[0]<=REG[0]<<0;
      10'h194: data = 32'h8fc20000; // 00400650: LW, REG[2]<=RAM[REG[30]+0];
      10'h195: data = 32'h00000000; // 00400654: SLL, REG[0]<=REG[0]<<0;
      10'h196: data = 32'h24420064; // 00400658: ADDIU, REG[2]<=REG[2]+100(=0x00000064);
      10'h197: data = 32'hafc20000; // 0040065c: SW, RAM[REG[30]+0]<=REG[2];
      10'h198: data = 32'h8fc20004; // 00400660: LW, REG[2]<=RAM[REG[30]+4];
      10'h199: data = 32'h00000000; // 00400664: SLL, REG[0]<=REG[0]<<0;
      10'h19a: data = 32'h24420001; // 00400668: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h19b: data = 32'hafc20004; // 0040066c: SW, RAM[REG[30]+4]<=REG[2];
      10'h19c: data = 32'h8fc20008; // 00400670: LW, REG[2]<=RAM[REG[30]+8];
      10'h19d: data = 32'h00000000; // 00400674: SLL, REG[0]<=REG[0]<<0;
      10'h19e: data = 32'h8c420000; // 00400678: LW, REG[2]<=RAM[REG[2]+0];
      10'h19f: data = 32'h00000000; // 0040067c: SLL, REG[0]<=REG[0]<<0;
      10'h1a0: data = 32'h2443ffd0; // 00400680: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h1a1: data = 32'h8fc20004; // 00400684: LW, REG[2]<=RAM[REG[30]+4];
      10'h1a2: data = 32'h00000000; // 00400688: SLL, REG[0]<=REG[0]<<0;
      10'h1a3: data = 32'h0043102b; // 0040068c: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h1a4: data = 32'h1440ffef; // 00400690: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h1a5: data = 32'h00000000; // 00400694: SLL, REG[0]<=REG[0]<<0;
      10'h1a6: data = 32'h8fc20008; // 00400698: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a7: data = 32'h00000000; // 0040069c: SLL, REG[0]<=REG[0]<<0;
      10'h1a8: data = 32'h24420004; // 004006a0: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h1a9: data = 32'hafc20008; // 004006a4: SW, RAM[REG[30]+8]<=REG[2];
      10'h1aa: data = 32'hafc00004; // 004006a8: SW, RAM[REG[30]+4]<=REG[0];
      10'h1ab: data = 32'h081001b5; // 004006ac: J, PC<=0x001001b5*4(=0x004006d4);
      10'h1ac: data = 32'h00000000; // 004006b0: SLL, REG[0]<=REG[0]<<0;
      10'h1ad: data = 32'h8fc20000; // 004006b4: LW, REG[2]<=RAM[REG[30]+0];
      10'h1ae: data = 32'h00000000; // 004006b8: SLL, REG[0]<=REG[0]<<0;
      10'h1af: data = 32'h2442000a; // 004006bc: ADDIU, REG[2]<=REG[2]+10(=0x0000000a);
      10'h1b0: data = 32'hafc20000; // 004006c0: SW, RAM[REG[30]+0]<=REG[2];
      10'h1b1: data = 32'h8fc20004; // 004006c4: LW, REG[2]<=RAM[REG[30]+4];
      10'h1b2: data = 32'h00000000; // 004006c8: SLL, REG[0]<=REG[0]<<0;
      10'h1b3: data = 32'h24420001; // 004006cc: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h1b4: data = 32'hafc20004; // 004006d0: SW, RAM[REG[30]+4]<=REG[2];
      10'h1b5: data = 32'h8fc20008; // 004006d4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b6: data = 32'h00000000; // 004006d8: SLL, REG[0]<=REG[0]<<0;
      10'h1b7: data = 32'h8c420000; // 004006dc: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b8: data = 32'h00000000; // 004006e0: SLL, REG[0]<=REG[0]<<0;
      10'h1b9: data = 32'h2443ffd0; // 004006e4: ADDIU, REG[3]<=REG[2]+65488(=0x0000ffd0);
      10'h1ba: data = 32'h8fc20004; // 004006e8: LW, REG[2]<=RAM[REG[30]+4];
      10'h1bb: data = 32'h00000000; // 004006ec: SLL, REG[0]<=REG[0]<<0;
      10'h1bc: data = 32'h0043102b; // 004006f0: SLTU, REG[2]<=(REG[2]<REG[3])?1:0;
      10'h1bd: data = 32'h1440ffef; // 004006f4: BNE, PC<=(REG[2] != REG[0])?PC+4+65519*4:PC+4;
      10'h1be: data = 32'h00000000; // 004006f8: SLL, REG[0]<=REG[0]<<0;
      10'h1bf: data = 32'h8fc20008; // 004006fc: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c0: data = 32'h00000000; // 00400700: SLL, REG[0]<=REG[0]<<0;
      10'h1c1: data = 32'h24420004; // 00400704: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h1c2: data = 32'hafc20008; // 00400708: SW, RAM[REG[30]+8]<=REG[2];
      10'h1c3: data = 32'h8fc20008; // 0040070c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c4: data = 32'h00000000; // 00400710: SLL, REG[0]<=REG[0]<<0;
      10'h1c5: data = 32'h8c430000; // 00400714: LW, REG[3]<=RAM[REG[2]+0];
      10'h1c6: data = 32'h8fc20000; // 00400718: LW, REG[2]<=RAM[REG[30]+0];
      10'h1c7: data = 32'h00000000; // 0040071c: SLL, REG[0]<=REG[0]<<0;
      10'h1c8: data = 32'h00621021; // 00400720: ADDU, REG[2]<=REG[3]+REG[2];
      10'h1c9: data = 32'h2442ffd0; // 00400724: ADDIU, REG[2]<=REG[2]+65488(=0x0000ffd0);
      10'h1ca: data = 32'hafc20000; // 00400728: SW, RAM[REG[30]+0]<=REG[2];
      10'h1cb: data = 32'h8fc20000; // 0040072c: LW, REG[2]<=RAM[REG[30]+0];
      10'h1cc: data = 32'h03c0e821; // 00400730: ADDU, REG[29]<=REG[30]+REG[0];
      10'h1cd: data = 32'h8fbe0010; // 00400734: LW, REG[30]<=RAM[REG[29]+16];
      10'h1ce: data = 32'h27bd0018; // 00400738: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h1cf: data = 32'h03e00008; // 0040073c: JR, PC<=REG[31];
      10'h1d0: data = 32'h00000000; // 00400740: SLL, REG[0]<=REG[0]<<0;
      10'h1d1: data = 32'h00000000; // 00400744: SLL, REG[0]<=REG[0]<<0;
      10'h1d2: data = 32'h00000000; // 00400748: SLL, REG[0]<=REG[0]<<0;
      10'h1d3: data = 32'h00000000; // 0040074c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
